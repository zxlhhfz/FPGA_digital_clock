module temp_humi_display(
    input PixelClk,
    input nRST,
    input [15:0] PixelCount,
    input [15:0] LineCount,
    input [31:0] TempHumi,
    input [15:0] temp, //温度值
    input [15:0] humi, //湿度值
    output reg [4:0] LCD_B,
    output reg [5:0] LCD_G,
    output reg [4:0] LCD_R
);

wire [0:39] wendu_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0600000200, 40'h0381800300, 40'h01C1FFFF00, 40'h00C1800300, 40'h00C1800300,
    40'h0001800300, 40'h0009800300, 40'h0009FFFF00, 40'h2009800300, 40'h1811800300, 40'h1C11800300, 40'h0E11800300, 40'h0E21800300,
    40'h0621800300, 40'h0421FFFF00, 40'h0061800300, 40'h0041800000, 40'h0040000000, 40'h00C40000C0, 40'h00C7FFFFE0, 40'h00861860C0,
    40'h01861860C0, 40'h01861860C0, 40'h23861860C0, 40'h1F061860C0, 40'h07061860C0, 40'h03061860C0, 40'h03061860C0, 40'h07061860C0,
    40'h07061860C0, 40'h07061860C8, 40'h07061860D8, 40'h07FFFFFFFC, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; //汉字“温”

wire [0:39] du_char [0:39] = '{
    40'h0000000000, 40'h0000300000, 40'h00001C0000, 40'h00000E0000, 40'h0000060020, 40'h0300060070, 40'h03FFFFFFF8, 40'h0380000000,
    40'h0380801000, 40'h0380E01C00, 40'h0380C01800, 40'h0380C01840, 40'h0380C018E0, 40'h03FFFFFFF0, 40'h0380C01800, 40'h0380C01800,
    40'h0300C01800, 40'h0300C01800, 40'h0300C01800, 40'h0300FFF800, 40'h0300C01800, 40'h0300000000, 40'h0300000600, 40'h030FFFFF00,
    40'h0300800E00, 40'h0600401C00, 40'h0600203800, 40'h0600307000, 40'h0600186000, 40'h04000CC000, 40'h0C00078000, 40'h0C00070000,
    40'h08000FC000, 40'h180038F800, 40'h1000E03F80, 40'h1007800FFC, 40'h203C0001E0, 40'h41C0000000, 40'h0000000000, 40'h0000000000
}; //汉字“度”

wire [0:39] du2_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h03E003C000, 40'h06203FF800, 40'h0430700E40,
    40'h0430E00340, 40'h0421C001C0, 40'h07638000C0, 40'h01C30000C0, 40'h0007000040, 40'h0007000040, 40'h0006000040, 40'h000E000040,
    40'h000E000000, 40'h000E000000, 40'h000E000000, 40'h000E000000, 40'h000E000000, 40'h000E000000, 40'h000E000000, 40'h000E000000,
    40'h0006000000, 40'h0007000000, 40'h0007000000, 40'h0003800040, 40'h0003800080, 40'h0001C00180, 40'h0000E00700, 40'h0000781C00,
    40'h00003FF800, 40'h000007C000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; //符号“℃”

wire [0:39] shidu_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0400000000, 40'h03018000C0, 40'h0381FFFFE0, 40'h01C1C000C0, 40'h00C1C000C0, 40'h00C1C000C0,
    40'h0001C000C0, 40'h0009C000C0, 40'h0009FFFFC0, 40'h2011C000C0, 40'h1811C000C0, 40'h0C11C000C0, 40'h0E21C000C0, 40'h0721C000C0,
    40'h0621FFFFC0, 40'h0241C000C0, 40'h00418C3000, 40'h00C00E3800, 40'h00800C3000, 40'h01880C3030, 40'h018C0C3038, 40'h03860C3070,
    40'h03030C30E0, 40'h3F038C30C0, 40'h0F038C3180, 40'h0701CC3300, 40'h0601CC3600, 40'h0600CC3400, 40'h06008C3800, 40'h0E000C3000,
    40'h0E000C3000, 40'h0E000C3010, 40'h0E000C3038, 40'h023FFFFFFC, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; //汉字“湿”

wire [0:39] baifenhao_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h01E0000400, 40'h07BC000E00,
    40'h1C07000C00, 40'h3C07801800, 40'h3807803000, 40'h7803C07000, 40'h7803C0E000, 40'h7803C1C000, 40'h7803C18000, 40'h7803C30000,
    40'h3807860000, 40'h3C078E0000, 40'h1C0F1C0000, 40'h071E180F00, 40'h00E03079E0, 40'h000061E070, 40'h0000C1C078, 40'h0001C3C038,
    40'h000383803C, 40'h000307803C, 40'h000607803C, 40'h000C07803C, 40'h001807803C, 40'h003803C03C, 40'h007001C078, 40'h006001E070,
    40'h00C00079E0, 40'h0080000F00, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; //符号“%”

wire [0:19] dian_char [0:39] = '{
    20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000,
    20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000,
    20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00600, 20'h00F00, 20'h00F00, 20'h00600, 20'h00000,
    20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000, 20'h00000
}; //符号“.”

wire [0:39] zero_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00007E0000, 40'h0007FFE000,    
    40'h001F007800, 40'h007C003E00, 40'h00F8001F00, 40'h01F0000F80, 40'h03F0000FC0, 40'h07E00007C0, 40'h07E00007E0, 40'h0FC00003E0,    
    40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0,    
    40'h0FC00003F0, 40'h0FC00003E0, 40'h07E00007E0, 40'h07E00007C0, 40'h03E0000FC0, 40'h01F0000F80, 40'h00F8001F00, 40'h007C003E00,    
    40'h001F00F800, 40'h0007FFE000, 40'h00007E0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] one_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000060000, 40'h00000E0000,
    40'h0000FE0000, 40'h007FFE0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000,
    40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000,
    40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00007F0000,
    40'h007FFFFF00, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};  

wire [0:39] two_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00007F0000, 40'h001F87F800,
    40'h0078003E00, 40'h01E0001F80, 40'h03C0000FC0, 40'h07C00007C0, 40'h07E00007C0, 40'h07F00007C0, 40'h03F00007C0, 40'h0000000FC0,
    40'h0000000F80, 40'h0000001F00, 40'h0000003C00, 40'h000000F800, 40'h000001E000, 40'h0000078000, 40'h00001E0000, 40'h0000780000,
    40'h0001E00000, 40'h0007800000, 40'h001E000000, 40'h0038000060, 40'h00E00000C0, 40'h03C00001C0, 40'h07000007C0, 40'h0FFFFFFFC0,
    40'h0FFFFFFF80, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; 

wire [0:39] three_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000FC0000, 40'h001F0FE000,
    40'h00F000F800, 40'h01E0003E00, 40'h03E0001F00, 40'h03F0001F80, 40'h03F0001F80, 40'h01E0001F80, 40'h0000001F00, 40'h0000001F00,
    40'h0000007C00, 40'h000001F000, 40'h00007F8000, 40'h0001FFC000, 40'h000000F800, 40'h0000001F00, 40'h0000000F80, 40'h00000007C0,
    40'h00000007E0, 40'h00000007E0, 40'h01C00007E0, 40'h07F00007E0, 40'h07F00007C0, 40'h07E0000F80, 40'h03E0001F00, 40'h01F0007C00,
    40'h003F07F000, 40'h0001FE0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] four_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000007800, 40'h000000F800,
    40'h000001F800, 40'h000003F800, 40'h00000EF800, 40'h00001CF800, 40'h000038F800, 40'h000060F800, 40'h0001C0F800, 40'h000380F800,
    40'h000700F800, 40'h000C00F800, 40'h003800F800, 40'h007000F800, 40'h00C000F800, 40'h018000F800, 40'h070000F800, 40'h0E0000F800,
    40'h1FFFFFFFF8, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000001F800,
    40'h0000FFFFF0, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; 

wire [0:39] five_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00FFFFFFC0,
    40'h00FFFFFF80, 40'h00E0000000, 40'h00C0000000, 40'h00C0000000, 40'h00C0000000, 40'h00C0000000, 40'h00C0000000, 40'h01C0000000,
    40'h01C07FC000, 40'h01C7FFF800, 40'h019C007E00, 40'h01F0001F80, 40'h01C0000FC0, 40'h00000007C0, 40'h00000007E0, 40'h00000003E0,
    40'h00000003E0, 40'h00000003E0, 40'h03E00003E0, 40'h07F00007C0, 40'h07E00007C0, 40'h07C0000F80, 40'h03C0001F00, 40'h00E0007E00,
    40'h003F87F000, 40'h0001FE0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; 

wire [0:39] six_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00000FC000, 40'h0001F8FC00,
    40'h000F001F00, 40'h003C001F80, 40'h0078001F80, 40'h01F0000E00, 40'h01E0000000, 40'h03E0000000, 40'h07C0000000, 40'h07C0000000,
    40'h0FC01F8000, 40'h0FC3FFFC00, 40'h0FCF803F00, 40'h0FDC000F80, 40'h0FF00007C0, 40'h0FE00003E0, 40'h0FC00003F0, 40'h0FC00001F0,
    40'h0FC00001F0, 40'h0FC00001F0, 40'h07C00003F0, 40'h07E00003E0, 40'h03E00003E0, 40'h01F00007C0, 40'h00FC000780, 40'h003E001E00,
    40'h000FE1F800, 40'h00007F0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] seven_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h01FFFFFFE0,
    40'h01FFFFFFC0, 40'h03E0000380, 40'h0380000700, 40'h0300000E00, 40'h0600001C00, 40'h0000003800, 40'h0000007000, 40'h000000E000,
    40'h000001C000, 40'h0000038000, 40'h0000078000, 40'h00000F0000, 40'h00001E0000, 40'h00003E0000, 40'h00003C0000, 40'h00007C0000,
    40'h0000F80000, 40'h0000F80000, 40'h0001F80000, 40'h0001F80000, 40'h0001F80000, 40'h0003F80000, 40'h0003F80000, 40'h0003F80000,
    40'h0003F80000, 40'h0000F00000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] eight_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000FF0000, 40'h001FC3F800,
    40'h00F8001E00, 40'h01E0000F80, 40'h03C00007C0, 40'h07800003C0, 40'h07800003E0, 40'h07C00003E0, 40'h07E00003C0, 40'h03F0000780,
    40'h01FE000F00, 40'h007FC03C00, 40'h001FFFE000, 40'h0007FFC000, 40'h003C1FF800, 40'h00F003FE00, 40'h03C0007F80, 40'h0780001FC0,
    40'h0F800007E0, 40'h0F000003E0, 40'h1F000001E0, 40'h1F000001E0, 40'h0F000003E0, 40'h07800003C0, 40'h03C0000780, 40'h00F0001E00,
    40'h003F83F800, 40'h0000FE0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] nine_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000FC0000, 40'h003F87E000,
    40'h00F8007C00, 40'h01E0001E00, 40'h07C0000F00, 40'h07C0000780, 40'h0F800007C0, 40'h0F800007E0, 40'h1F800003E0, 40'h1F800003E0,
    40'h0F800003E0, 40'h0F800007F0, 40'h0FC0000FF0, 40'h07E0001BF0, 40'h03F00073F0, 40'h01FC03C7E0, 40'h003FFF07E0, 40'h00000007E0,
    40'h00000007C0, 40'h0000000FC0, 40'h0000000F80, 40'h0000001F00, 40'h00E0001E00, 40'h01F0003C00, 40'h03F800F800, 40'h01F803E000,
    40'h007E3F8000, 40'h0007F00000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

    wire [3:0] temp_first;
    wire [3:0] temp_second;
    wire [3:0] temp_third;
    wire [3:0] temp_fourth;
    wire [3:0] humi_first;
    wire [3:0] humi_second;
    wire [3:0] humi_third;
    wire [3:0] humi_fourth;
    
    assign temp_first = TempHumi[31:24] / 10;
    assign temp_second = TempHumi[31:24] % 10;
    assign temp_third = TempHumi[23:16] / 10;
    assign temp_fourth = TempHumi[23:16] % 10;
    assign humi_first = TempHumi[15:8] / 10;
    assign humi_second = TempHumi[15:8] % 10;
    assign humi_third = TempHumi[7:0] / 10;
    assign humi_fourth = TempHumi[7:0] % 10;

    localparam DISPLAY_Y1_START = 180;
    localparam DISPLAY_Y1_END = 220;
    localparam DISPLAY_Y2_START = 230;
    localparam DISPLAY_Y2_END = 270;

    function automatic get_digit_pixel;
        input [3:0] digit;
        input [15:0] x_pos;
        input [15:0] y_pos;
        reg pixel;
        begin
            case(digit)
                4'd0: pixel = zero_char[y_pos][x_pos];
                4'd1: pixel = one_char[y_pos][x_pos];
                4'd2: pixel = two_char[y_pos][x_pos];
                4'd3: pixel = three_char[y_pos][x_pos];
                4'd4: pixel = four_char[y_pos][x_pos];
                4'd5: pixel = five_char[y_pos][x_pos];
                4'd6: pixel = six_char[y_pos][x_pos];
                4'd7: pixel = seven_char[y_pos][x_pos];
                4'd8: pixel = eight_char[y_pos][x_pos];
                4'd9: pixel = nine_char[y_pos][x_pos];
                default: pixel = 1'b0;
            endcase
            get_digit_pixel = pixel;
        end
    endfunction

    always @(posedge PixelClk or negedge nRST) begin
        if(!nRST) begin
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
        end
        else if(LineCount >= DISPLAY_Y1_START && LineCount < DISPLAY_Y1_END) begin
            // 计算相对位置
            integer x_pos = PixelCount - 190; // 基准偏移
            integer y_pos = LineCount - DISPLAY_Y1_START;
            
            // 默认背景色
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
            
            // 汉字"温度"显示
            if(PixelCount >= 190 && PixelCount < 230) begin
                if(wendu_char[y_pos][x_pos]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
            else if(PixelCount >= 230 && PixelCount < 270) begin
                if(du_char[y_pos][x_pos-40]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
           
            // 温度整数显示
            else if(PixelCount >= 280 && PixelCount < 320) begin
                if(get_digit_pixel(temp_first, x_pos-90, y_pos))
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end
            else if(PixelCount >= 320 && PixelCount < 360) begin
                if(get_digit_pixel(temp_second, x_pos-130, y_pos))
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end
            
 //           点号显示
//            else if(PixelCount >= 360 && PixelCount < 380) begin
//                integer colon_x = PixelCount - 360;
//                if(dian_char[y_pos][colon_x])
//                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
//            end
//            
//             温度小数显示
//            else if(PixelCount >= 380 && PixelCount < 420) begin
//                if(get_digit_pixel(temp_third, x_pos-190, y_pos))
//                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
//            end
//            else if(PixelCount >= 420 && PixelCount < 460) begin
//                if(get_digit_pixel(temp_fourth, x_pos-230, y_pos))
//                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
//            end

             // 摄氏度显示
            else if(PixelCount >= 360 && PixelCount < 400) begin
                integer colon_x = PixelCount - 360;
                if(du2_char[y_pos][colon_x])
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end 
          
        end
        else if(LineCount >= DISPLAY_Y2_START && LineCount < DISPLAY_Y2_END) begin
            // 计算相对位置
            integer x_pos = PixelCount - 190; // 基准偏移
            integer y_pos = LineCount - DISPLAY_Y2_START;
            
            // 默认背景色
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
            
            // 汉字"湿度"显示
            if(PixelCount >= 190 && PixelCount < 230) begin
                if(shidu_char[y_pos][x_pos]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
            else if(PixelCount >= 230 && PixelCount < 270) begin
                if(du_char[y_pos][x_pos-40]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
           
            // 温度整数显示
            else if(PixelCount >= 280 && PixelCount < 320) begin
                if(get_digit_pixel(humi_first, x_pos-90, y_pos))
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end
            else if(PixelCount >= 320 && PixelCount < 360) begin
                if(get_digit_pixel(humi_second, x_pos-130, y_pos))
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end
            
//             点号显示
//            else if(PixelCount >= 360 && PixelCount < 380) begin
//                integer colon_x = PixelCount - 360;
//                if(dian_char[y_pos][colon_x])
//                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
//            end
//            
//             温度小数显示
//            else if(PixelCount >= 380 && PixelCount < 420) begin
//                if(get_digit_pixel(humi_third, x_pos-190, y_pos))
//                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
//            end
//            else if(PixelCount >= 420 && PixelCount < 460) begin
//                if(get_digit_pixel(humi_fourth, x_pos-230, y_pos))
//                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
//            end

             // 百分号显示
            else if(PixelCount >= 360 && PixelCount < 400) begin
                integer colon_x = PixelCount - 360;
                if(baifenhao_char[y_pos][colon_x])
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end 
          
        end
        else begin
            // 非显示区域
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
        end
    end    

endmodule