module alarm_hourly_display(
    input PixelClk,
    input nRST,
    input [15:0] PixelCount,
    input [15:0] LineCount,
    input [5:0] hour_decimal,
    input [5:0] alarm_hourly_en,
    output reg [4:0] LCD_B,
    output reg [5:0] LCD_G,
    output reg [4:0] LCD_R
);

    // 显示区域参数
    localparam DISPLAY_X_START = 190;
    localparam DISPLAY_X_END = 400;
    localparam DISPLAY_Y_START = 280;
    localparam DISPLAY_Y_END = 320;

wire [0:39] shi_char [0:39] = '{
    40'h0000000000, 40'h0000000800, 40'h0000000E00, 40'h0000000E00, 40'h0000000C00, 40'h0000000C00, 40'h180C000C00, 40'h1FFF000C00,
    40'h0C0E000C00, 40'h0C0C000C20, 40'h0C0C000C70, 40'h0C0DFFFFF8, 40'h0C0C000C00, 40'h0C0C000C00, 40'h0C0C000C00, 40'h0C0C000C00,
    40'h0C0C200C00, 40'h0FFC300C00, 40'h0C0C180C00, 40'h0C0C1C0C00, 40'h0C0C0E0C00, 40'h0C0C0E0C00, 40'h0C0C060C00, 40'h0C0C060C00,
    40'h0C0C060C00, 40'h0C0C000C00, 40'h0C0C000C00, 40'h0C0C000C00, 40'h0C0C000C00, 40'h0FFC000C00, 40'h0C0C000C00, 40'h0C0E000C00,
    40'h1C08000C00, 40'h1800000C00, 40'h000003FC00, 40'h0000007C00, 40'h0000003800, 40'h0000001000, 40'h0000000000, 40'h0000000000
}; //汉字“时”

wire [0:39] bao_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0040000000, 40'h0070300100, 40'h00603FFF80, 40'h0060380380, 40'h0060380300, 40'h0060380300,
    40'h0060380300, 40'h0060380300, 40'h0063380300, 40'h3FFFB80300, 40'h0060784700, 40'h0060383E00, 40'h0060381E00, 40'h0060380800,
    40'h00603800C0, 40'h0061BFFFE0, 40'h00663901C0, 40'h0078390180, 40'h01E0390180, 40'h0FE0388300, 40'h3E60388300, 40'h186038C600,
    40'h1060384600, 40'h0060386C00, 40'h0060383C00, 40'h0060381800, 40'h0060383C00, 40'h0060387E00, 40'h006038E700, 40'h006038C3C0,
    40'h00603901F0, 40'h00603E00FC, 40'h1FE03C0030, 40'h07E0380000, 40'h01C0300000, 40'h0080000000, 40'h0000000000, 40'h0000000000
}; //汉字“报”

wire [0:39] zhong_image [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h3C0000003C, 40'h6600000066, 40'h52000000DA, 40'h5BFFFFFF32, 40'h4BFFFFFFA2, 40'h67FFFFFFEC,
    40'h3C00000070, 40'h1C00000070, 40'h1C00100070, 40'h1C00300070, 40'h1C00100070, 40'h1C00100070, 40'h1C00100070, 40'h1C0010C070,
    40'h1C0011FC70, 40'h1C00178070, 40'h1C003E0070, 40'h1C003C0070, 40'h1C00380070, 40'h1C00380070, 40'h1C00000070, 40'h1C00000070,
    40'h1C00000070, 40'h1C00000070, 40'h1C00000070, 40'h1C00000070, 40'h1C00000070, 40'h1C00000070, 40'h1C00000070, 40'h1E000000F0,
    40'h0F000001E0, 40'h07FFFFFFC0, 40'h01FFFFFF00, 40'h01FFFFFF00, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; //闹钟图形

wire [0:39] zero_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00007E0000, 40'h0007FFE000,    
    40'h001F007800, 40'h007C003E00, 40'h00F8001F00, 40'h01F0000F80, 40'h03F0000FC0, 40'h07E00007C0, 40'h07E00007E0, 40'h0FC00003E0,    
    40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0, 40'h0FC00003F0,    
    40'h0FC00003F0, 40'h0FC00003E0, 40'h07E00007E0, 40'h07E00007C0, 40'h03E0000FC0, 40'h01F0000F80, 40'h00F8001F00, 40'h007C003E00,    
    40'h001F00F800, 40'h0007FFE000, 40'h00007E0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] one_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000060000, 40'h00000E0000,
    40'h0000FE0000, 40'h007FFE0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000,
    40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000,
    40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00003E0000, 40'h00007F0000,
    40'h007FFFFF00, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};  

wire [0:39] two_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00007F0000, 40'h001F87F800,
    40'h0078003E00, 40'h01E0001F80, 40'h03C0000FC0, 40'h07C00007C0, 40'h07E00007C0, 40'h07F00007C0, 40'h03F00007C0, 40'h0000000FC0,
    40'h0000000F80, 40'h0000001F00, 40'h0000003C00, 40'h000000F800, 40'h000001E000, 40'h0000078000, 40'h00001E0000, 40'h0000780000,
    40'h0001E00000, 40'h0007800000, 40'h001E000000, 40'h0038000060, 40'h00E00000C0, 40'h03C00001C0, 40'h07000007C0, 40'h0FFFFFFFC0,
    40'h0FFFFFFF80, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; 

wire [0:39] three_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000FC0000, 40'h001F0FE000,
    40'h00F000F800, 40'h01E0003E00, 40'h03E0001F00, 40'h03F0001F80, 40'h03F0001F80, 40'h01E0001F80, 40'h0000001F00, 40'h0000001F00,
    40'h0000007C00, 40'h000001F000, 40'h00007F8000, 40'h0001FFC000, 40'h000000F800, 40'h0000001F00, 40'h0000000F80, 40'h00000007C0,
    40'h00000007E0, 40'h00000007E0, 40'h01C00007E0, 40'h07F00007E0, 40'h07F00007C0, 40'h07E0000F80, 40'h03E0001F00, 40'h01F0007C00,
    40'h003F07F000, 40'h0001FE0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] four_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000007800, 40'h000000F800,
    40'h000001F800, 40'h000003F800, 40'h00000EF800, 40'h00001CF800, 40'h000038F800, 40'h000060F800, 40'h0001C0F800, 40'h000380F800,
    40'h000700F800, 40'h000C00F800, 40'h003800F800, 40'h007000F800, 40'h00C000F800, 40'h018000F800, 40'h070000F800, 40'h0E0000F800,
    40'h1FFFFFFFF8, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000000F800, 40'h000001F800,
    40'h0000FFFFF0, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; 

wire [0:39] five_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00FFFFFFC0,
    40'h00FFFFFF80, 40'h00E0000000, 40'h00C0000000, 40'h00C0000000, 40'h00C0000000, 40'h00C0000000, 40'h00C0000000, 40'h01C0000000,
    40'h01C07FC000, 40'h01C7FFF800, 40'h019C007E00, 40'h01F0001F80, 40'h01C0000FC0, 40'h00000007C0, 40'h00000007E0, 40'h00000003E0,
    40'h00000003E0, 40'h00000003E0, 40'h03E00003E0, 40'h07F00007C0, 40'h07E00007C0, 40'h07C0000F80, 40'h03C0001F00, 40'h00E0007E00,
    40'h003F87F000, 40'h0001FE0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
}; 

wire [0:39] six_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h00000FC000, 40'h0001F8FC00,
    40'h000F001F00, 40'h003C001F80, 40'h0078001F80, 40'h01F0000E00, 40'h01E0000000, 40'h03E0000000, 40'h07C0000000, 40'h07C0000000,
    40'h0FC01F8000, 40'h0FC3FFFC00, 40'h0FCF803F00, 40'h0FDC000F80, 40'h0FF00007C0, 40'h0FE00003E0, 40'h0FC00003F0, 40'h0FC00001F0,
    40'h0FC00001F0, 40'h0FC00001F0, 40'h07C00003F0, 40'h07E00003E0, 40'h03E00003E0, 40'h01F00007C0, 40'h00FC000780, 40'h003E001E00,
    40'h000FE1F800, 40'h00007F0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] seven_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h01FFFFFFE0,
    40'h01FFFFFFC0, 40'h03E0000380, 40'h0380000700, 40'h0300000E00, 40'h0600001C00, 40'h0000003800, 40'h0000007000, 40'h000000E000,
    40'h000001C000, 40'h0000038000, 40'h0000078000, 40'h00000F0000, 40'h00001E0000, 40'h00003E0000, 40'h00003C0000, 40'h00007C0000,
    40'h0000F80000, 40'h0000F80000, 40'h0001F80000, 40'h0001F80000, 40'h0001F80000, 40'h0003F80000, 40'h0003F80000, 40'h0003F80000,
    40'h0003F80000, 40'h0000F00000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] eight_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000FF0000, 40'h001FC3F800,
    40'h00F8001E00, 40'h01E0000F80, 40'h03C00007C0, 40'h07800003C0, 40'h07800003E0, 40'h07C00003E0, 40'h07E00003C0, 40'h03F0000780,
    40'h01FE000F00, 40'h007FC03C00, 40'h001FFFE000, 40'h0007FFC000, 40'h003C1FF800, 40'h00F003FE00, 40'h03C0007F80, 40'h0780001FC0,
    40'h0F800007E0, 40'h0F000003E0, 40'h1F000001E0, 40'h1F000001E0, 40'h0F000003E0, 40'h07800003C0, 40'h03C0000780, 40'h00F0001E00,
    40'h003F83F800, 40'h0000FE0000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};

wire [0:39] nine_char [0:39] = '{
    40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000FC0000, 40'h003F87E000,
    40'h00F8007C00, 40'h01E0001E00, 40'h07C0000F00, 40'h07C0000780, 40'h0F800007C0, 40'h0F800007E0, 40'h1F800003E0, 40'h1F800003E0,
    40'h0F800003E0, 40'h0F800007F0, 40'h0FC0000FF0, 40'h07E0001BF0, 40'h03F00073F0, 40'h01FC03C7E0, 40'h003FFF07E0, 40'h00000007E0,
    40'h00000007C0, 40'h0000000FC0, 40'h0000000F80, 40'h0000001F00, 40'h00E0001E00, 40'h01F0003C00, 40'h03F800F800, 40'h01F803E000,
    40'h007E3F8000, 40'h0007F00000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000, 40'h0000000000
};
    
    // 数字分解
    wire [3:0] hour_first = hour_decimal / 10;
    wire [3:0] hour_second = hour_decimal % 10;

    // 闹钟激活标志
    wire alarm_active = (alarm_hourly_en > 0) && ((alarm_hourly_en - 1'd1) % 2 == 0) && 
                       (alarm_hourly_en < 6'd1 + hour_decimal * 2);

    // 显示数字的函数
    function automatic [15:0] get_digit_pixel;
        input [3:0] digit;
        input [15:0] x_pos;
        input [15:0] y_pos;
        begin
            case(digit)
                4'd0: get_digit_pixel = zero_char[y_pos][x_pos];
                4'd1: get_digit_pixel = one_char[y_pos][x_pos];
                4'd2: get_digit_pixel = two_char[y_pos][x_pos];
                4'd3: get_digit_pixel = three_char[y_pos][x_pos];
                4'd4: get_digit_pixel = four_char[y_pos][x_pos];
                4'd5: get_digit_pixel = five_char[y_pos][x_pos];
                4'd6: get_digit_pixel = six_char[y_pos][x_pos];
                4'd7: get_digit_pixel = seven_char[y_pos][x_pos];
                4'd8: get_digit_pixel = eight_char[y_pos][x_pos];
                4'd9: get_digit_pixel = nine_char[y_pos][x_pos];
                default: get_digit_pixel = 1'b0;
            endcase
        end
    endfunction

    // 主显示逻辑
    always @(posedge PixelClk or negedge nRST) begin
        if(!nRST) begin
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
        end
        else if(LineCount >= DISPLAY_Y_START && LineCount < DISPLAY_Y_END) begin
            // 计算相对位置
            integer x_pos = PixelCount - DISPLAY_X_START;
            integer y_pos = LineCount - DISPLAY_Y_START;
            
            // 默认背景色
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
            
            // "报"字显示区域 (190-230)
            if(PixelCount >= 190 && PixelCount < 230) begin
                if(bao_char[y_pos][x_pos]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
            // "时"字显示区域 (230-270)
            else if(PixelCount >= 230 && PixelCount < 270) begin
                if(shi_char[y_pos][x_pos-40]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
            // 闹钟图标显示区域 (280-320)
            else if(PixelCount >= 280 && PixelCount < 320) begin
                if(alarm_active && zhong_image[y_pos][x_pos-90]) 
                    {LCD_R, LCD_G, LCD_B} <= {5'b00000, 6'b000000, 5'b00000};
            end
            // 小时十位数显示区域 (320-360)
            else if(PixelCount >= 320 && PixelCount < 360) begin
                if(alarm_active && get_digit_pixel(hour_first, x_pos-130, y_pos))
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end
            // 小时个位数显示区域 (360-400)
            else if(PixelCount >= 360 && PixelCount < 400) begin
                if(alarm_active && get_digit_pixel(hour_second, x_pos-170, y_pos))
                    {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b000000, 5'b00000};
            end
        end
        else begin
            // 非显示区域
            {LCD_R, LCD_G, LCD_B} <= {5'b11111, 6'b111111, 5'b11111};
        end
    end
endmodule