module clock_image_display(
    input PixelClk,
    input nRST,
    input [15:0] PixelCount,
    input [15:0] LineCount,
    output reg [4:0] LCD_B,
    output reg [5:0] LCD_G,
    output reg [4:0] LCD_R,

    input   [5:0]   hour_decimal,
    input   [5:0]   minute_decimal,
    input   [5:0]   second_decimal
);

wire [0:79] hour_000 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h0000000001c000000000, 80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000,
    80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000,
    80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000,
    80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003e000000000,
    80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000001c000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_030 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000780000000, 80'h00000000000780000000,
    80'h00000000000fc0000000, 80'h00000000000fc0000000, 80'h00000000001f80000000, 80'h00000000001f00000000,
    80'h00000000003f00000000, 80'h00000000007e00000000, 80'h00000000007e00000000, 80'h0000000000fc00000000,
    80'h0000000000f800000000, 80'h0000000001f800000000, 80'h0000000001f000000000, 80'h0000000003f000000000,
    80'h0000000003e000000000, 80'h0000000003e000000000, 80'h0000000003c000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_060 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000018000000,
    80'h0000000000007c000000, 80'h000000000001fe000000, 80'h000000000003fc000000, 80'h00000000000ffc000000,
    80'h00000000003ff0000000, 80'h0000000000ffc0000000, 80'h0000000001ff80000000, 80'h0000000003fe00000000,
    80'h0000000007f800000000, 80'h0000000007e000000000, 80'h0000000003c000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_090 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003fffe000000, 80'h0000000007ffff000000,
    80'h0000000007ffff000000, 80'h0000000007ffff000000, 80'h0000000003fffe000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_120 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000078000000000, 80'h0000000007e000000000,
    80'h0000000007f800000000, 80'h0000000007fe00000000, 80'h0000000003ff00000000, 80'h0000000000ffc0000000,
    80'h00000000003ff0000000, 80'h00000000000ffc000000, 80'h000000000007fc000000, 80'h000000000001fc000000,
    80'h0000000000007c000000, 80'h00000000000030000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_150 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000030000000000, 80'h00000000078000000000, 80'h0000000007c000000000,
    80'h0000000007e000000000, 80'h0000000007e000000000, 80'h0000000003f000000000, 80'h0000000001f000000000,
    80'h0000000001f800000000, 80'h0000000000f800000000, 80'h0000000000fc00000000, 80'h00000000007e00000000,
    80'h00000000007e00000000, 80'h00000000003f00000000, 80'h00000000001f00000000, 80'h00000000001f80000000,
    80'h00000000000f80000000, 80'h00000000000f00000000, 80'h00000000000200000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_180 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000038000000000, 80'h0000000007c000000000, 80'h0000000007c000000000,
    80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000,
    80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000,
    80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000,
    80'h0000000007c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000, 80'h00000000038000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_210 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h0000000003c000000000, 80'h0000000007c000000000, 80'h0000000007c000000000,
    80'h000000000fc000000000, 80'h000000000f8000000000, 80'h000000001f8000000000, 80'h000000001f0000000000,
    80'h000000003f0000000000, 80'h000000007e0000000000, 80'h000000007e0000000000, 80'h00000000fc0000000000,
    80'h00000000f80000000000, 80'h00000001f80000000000, 80'h00000003f00000000000, 80'h00000003f00000000000,
    80'h00000001e00000000000, 80'h00000001e00000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_240 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h0000000003c000000000, 80'h0000000007e000000000, 80'h000000001fe000000000,
    80'h000000007fc000000000, 80'h00000001ff8000000000, 80'h00000003ff0000000000, 80'h0000000ffc0000000000,
    80'h0000003ff00000000000, 80'h0000003fc00000000000, 80'h0000007f800000000000, 80'h0000003e000000000000,
    80'h00000018000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_270 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h0000007fffc000000000, 80'h000000ffffe000000000, 80'h000000ffffe000000000,
    80'h000000ffffe000000000, 80'h0000007fffc000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_300 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000c000000000000, 80'h0000003e000000000000,
    80'h0000003f800000000000, 80'h0000003fe00000000000, 80'h0000003ff00000000000, 80'h0000000ffc0000000000,
    80'h00000003ff0000000000, 80'h00000000ffc000000000, 80'h000000007fe000000000, 80'h000000001fe000000000,
    80'h0000000007e000000000, 80'h0000000001e000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] hour_330 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000400000000000, 80'h00000000f00000000000, 80'h00000001f00000000000,
    80'h00000001f80000000000, 80'h00000000f80000000000, 80'h00000000fc0000000000, 80'h000000007e0000000000,
    80'h000000007e0000000000, 80'h000000003f0000000000, 80'h000000001f0000000000, 80'h000000001f8000000000,
    80'h000000000f8000000000, 80'h000000000fc000000000, 80'h0000000007e000000000, 80'h0000000007e000000000,
    80'h0000000003e000000000, 80'h0000000001e000000000, 80'h0000000000c000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};



wire [0:79] second_000 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_006 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000800000000, 80'h00000000000800000000, 80'h00000000001800000000, 80'h00000000001800000000,
    80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001000000000,
    80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000003000000000,
    80'h00000000003000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000002000000000, 80'h00000000006000000000, 80'h00000000006000000000, 80'h00000000004000000000,
    80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000004000000000,
    80'h00000000004000000000, 80'h00000000004000000000, 80'h0000000000c000000000, 80'h0000000000c000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_012 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000100000000, 80'h00000000000100000000, 80'h00000000000100000000,
    80'h00000000000100000000, 80'h00000000000300000000, 80'h00000000000200000000, 80'h00000000000200000000,
    80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000600000000, 80'h00000000000400000000,
    80'h00000000000400000000, 80'h00000000000400000000, 80'h00000000000c00000000, 80'h00000000000800000000,
    80'h00000000000800000000, 80'h00000000000800000000, 80'h00000000000800000000, 80'h00000000001800000000,
    80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001000000000,
    80'h00000000003000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000006000000000, 80'h00000000006000000000, 80'h00000000004000000000, 80'h00000000004000000000,
    80'h00000000004000000000, 80'h0000000000c000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_018 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000010000000, 80'h00000000000030000000,
    80'h00000000000020000000, 80'h00000000000020000000, 80'h00000000000060000000, 80'h00000000000040000000,
    80'h00000000000040000000, 80'h00000000000040000000, 80'h00000000000080000000, 80'h00000000000080000000,
    80'h00000000000080000000, 80'h00000000000100000000, 80'h00000000000100000000, 80'h00000000000100000000,
    80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000600000000,
    80'h00000000000400000000, 80'h00000000000400000000, 80'h00000000000c00000000, 80'h00000000000800000000,
    80'h00000000000800000000, 80'h00000000001800000000, 80'h00000000001000000000, 80'h00000000001000000000,
    80'h00000000003000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000006000000000,
    80'h00000000004000000000, 80'h00000000004000000000, 80'h0000000000c000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_024 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000002000000,
    80'h00000000000002000000, 80'h00000000000006000000, 80'h00000000000004000000, 80'h00000000000004000000,
    80'h00000000000008000000, 80'h00000000000008000000, 80'h00000000000018000000, 80'h00000000000010000000,
    80'h00000000000030000000, 80'h00000000000020000000, 80'h00000000000060000000, 80'h00000000000040000000,
    80'h00000000000040000000, 80'h00000000000080000000, 80'h00000000000080000000, 80'h00000000000180000000,
    80'h00000000000100000000, 80'h00000000000300000000, 80'h00000000000200000000, 80'h00000000000600000000,
    80'h00000000000400000000, 80'h00000000000400000000, 80'h00000000000800000000, 80'h00000000000800000000,
    80'h00000000001800000000, 80'h00000000001000000000, 80'h00000000003000000000, 80'h00000000002000000000,
    80'h00000000006000000000, 80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_030 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000600000, 80'h00000000000000400000, 80'h00000000000000c00000,
    80'h00000000000000800000, 80'h00000000000001800000, 80'h00000000000001000000, 80'h00000000000002000000,
    80'h00000000000006000000, 80'h00000000000004000000, 80'h0000000000000c000000, 80'h00000000000008000000,
    80'h00000000000018000000, 80'h00000000000010000000, 80'h00000000000020000000, 80'h00000000000060000000,
    80'h00000000000040000000, 80'h000000000000c0000000, 80'h00000000000080000000, 80'h00000000000100000000,
    80'h00000000000100000000, 80'h00000000000200000000, 80'h00000000000600000000, 80'h00000000000400000000,
    80'h00000000000c00000000, 80'h00000000000800000000, 80'h00000000001000000000, 80'h00000000003000000000,
    80'h00000000002000000000, 80'h00000000006000000000, 80'h00000000004000000000, 80'h0000000000c000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_036 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000040000,
    80'h00000000000000080000, 80'h00000000000000180000, 80'h00000000000000300000, 80'h00000000000000200000,
    80'h00000000000000400000, 80'h00000000000000c00000, 80'h00000000000001800000, 80'h00000000000001000000,
    80'h00000000000003000000, 80'h00000000000006000000, 80'h00000000000004000000, 80'h00000000000008000000,
    80'h00000000000018000000, 80'h00000000000030000000, 80'h00000000000020000000, 80'h00000000000040000000,
    80'h000000000000c0000000, 80'h00000000000080000000, 80'h00000000000100000000, 80'h00000000000300000000,
    80'h00000000000600000000, 80'h00000000000400000000, 80'h00000000000800000000, 80'h00000000001800000000,
    80'h00000000003000000000, 80'h00000000002000000000, 80'h00000000004000000000, 80'h0000000000c000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_042 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000010000, 80'h00000000000000030000,
    80'h00000000000000060000, 80'h000000000000000c0000, 80'h00000000000000180000, 80'h00000000000000300000,
    80'h00000000000000600000, 80'h00000000000000400000, 80'h00000000000000800000, 80'h00000000000001000000,
    80'h00000000000002000000, 80'h00000000000006000000, 80'h0000000000000c000000, 80'h00000000000018000000,
    80'h00000000000030000000, 80'h00000000000060000000, 80'h000000000000c0000000, 80'h00000000000080000000,
    80'h00000000000100000000, 80'h00000000000200000000, 80'h00000000000400000000, 80'h00000000000c00000000,
    80'h00000000001800000000, 80'h00000000003000000000, 80'h00000000006000000000, 80'h0000000000c000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_048 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000002000, 80'h00000000000000006000, 80'h0000000000000000c000, 80'h00000000000000010000,
    80'h00000000000000020000, 80'h000000000000000c0000, 80'h00000000000000180000, 80'h00000000000000300000,
    80'h00000000000000600000, 80'h00000000000000c00000, 80'h00000000000001800000, 80'h00000000000003000000,
    80'h00000000000004000000, 80'h00000000000008000000, 80'h00000000000030000000, 80'h00000000000060000000,
    80'h000000000000c0000000, 80'h00000000000180000000, 80'h00000000000300000000, 80'h00000000000600000000,
    80'h00000000000c00000000, 80'h00000000001000000000, 80'h00000000002000000000, 80'h0000000000c000000000,
    80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_054 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000c00,
    80'h00000000000000001800, 80'h00000000000000006000, 80'h0000000000000000c000, 80'h00000000000000018000,
    80'h00000000000000060000, 80'h000000000000000c0000, 80'h00000000000000300000, 80'h00000000000000600000,
    80'h00000000000000c00000, 80'h00000000000003000000, 80'h00000000000006000000, 80'h0000000000000c000000,
    80'h00000000000030000000, 80'h00000000000060000000, 80'h00000000000180000000, 80'h00000000000300000000,
    80'h00000000000600000000, 80'h00000000001800000000, 80'h00000000003000000000, 80'h00000000006000000000,
    80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_060 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000200, 80'h00000000000000000e00,
    80'h00000000000000001800, 80'h00000000000000006000, 80'h0000000000000001c000, 80'h00000000000000070000,
    80'h000000000000000c0000, 80'h00000000000000300000, 80'h00000000000000e00000, 80'h00000000000001800000,
    80'h00000000000006000000, 80'h00000000000018000000, 80'h00000000000070000000, 80'h000000000000c0000000,
    80'h00000000000300000000, 80'h00000000000e00000000, 80'h00000000003800000000, 80'h00000000006000000000,
    80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_066 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000080, 80'h00000000000000000380, 80'h00000000000000000e00,
    80'h00000000000000003800, 80'h0000000000000001c000, 80'h00000000000000070000, 80'h000000000000001c0000,
    80'h00000000000000700000, 80'h00000000000003800000, 80'h0000000000000e000000, 80'h00000000000038000000,
    80'h000000000000e0000000, 80'h00000000000700000000, 80'h00000000001c00000000, 80'h00000000007000000000,
    80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_072 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h000000000000000000c0, 80'h00000000000000000780, 80'h00000000000000003c00,
    80'h0000000000000001e000, 80'h000000000000000f0000, 80'h00000000000000700000, 80'h00000000000003800000,
    80'h0000000000003c000000, 80'h000000000001e0000000, 80'h00000000000f00000000, 80'h00000000007800000000,
    80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_078 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h000000000000000003e0, 80'h00000000000000007e00, 80'h0000000000000007c000,
    80'h00000000000000fc0000, 80'h0000000000001f800000, 80'h000000000001f0000000, 80'h00000000003f00000000,
    80'h0000000001e000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_084 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h000000000000000000f0, 80'h0000000000000001ffc0, 80'h00000000000007ff8000, 80'h00000000000ffe000000,
    80'h0000000001fc00000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_090 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h0000000001fffffffff0, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_096 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h0000000001fc00000000, 80'h00000000000ffe000000, 80'h00000000000007ff8000, 80'h0000000000000001ffc0,
    80'h000000000000000000f0, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_102 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h0000000001e000000000, 80'h00000000003f00000000, 80'h000000000003f0000000, 80'h0000000000001f800000,
    80'h00000000000000fc0000, 80'h0000000000000007c000, 80'h00000000000000007e00, 80'h000000000000000003e0,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_108 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h0000000001c000000000, 80'h00000000007800000000, 80'h00000000000f00000000, 80'h000000000001e0000000,
    80'h0000000000003c000000, 80'h00000000000007800000, 80'h00000000000000f00000, 80'h000000000000000e0000,
    80'h0000000000000001c000, 80'h00000000000000003c00, 80'h00000000000000000780, 80'h000000000000000000c0,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_114 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000018000000000, 80'h00000000007000000000, 80'h00000000001c00000000, 80'h00000000000700000000,
    80'h000000000001c0000000, 80'h00000000000038000000, 80'h0000000000000e000000, 80'h00000000000003800000,
    80'h00000000000000e00000, 80'h000000000000001c0000, 80'h00000000000000070000, 80'h0000000000000001c000,
    80'h00000000000000007000, 80'h00000000000000000e00, 80'h00000000000000000380, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_120 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000018000000000, 80'h0000000000e000000000, 80'h00000000003800000000, 80'h00000000000c00000000,
    80'h00000000000300000000, 80'h000000000001c0000000, 80'h00000000000060000000, 80'h00000000000018000000,
    80'h00000000000006000000, 80'h00000000000003800000, 80'h00000000000000c00000, 80'h00000000000000300000,
    80'h000000000000001c0000, 80'h00000000000000070000, 80'h00000000000000018000, 80'h00000000000000006000,
    80'h00000000000000003800, 80'h00000000000000000e00, 80'h00000000000000000200, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_126 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000018000000000, 80'h0000000000c000000000, 80'h00000000003000000000, 80'h00000000001800000000,
    80'h00000000000c00000000, 80'h00000000000300000000, 80'h00000000000180000000, 80'h000000000000c0000000,
    80'h00000000000030000000, 80'h00000000000018000000, 80'h00000000000006000000, 80'h00000000000003000000,
    80'h00000000000001800000, 80'h00000000000000600000, 80'h00000000000000300000, 80'h000000000000001c0000,
    80'h00000000000000060000, 80'h00000000000000030000, 80'h0000000000000000c000, 80'h00000000000000006000,
    80'h00000000000000003000, 80'h00000000000000000800, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_132 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000018000000000, 80'h0000000000c000000000, 80'h00000000006000000000, 80'h00000000003000000000,
    80'h00000000001800000000, 80'h00000000000c00000000, 80'h00000000000200000000, 80'h00000000000100000000,
    80'h000000000000c0000000, 80'h00000000000060000000, 80'h00000000000030000000, 80'h00000000000018000000,
    80'h0000000000000c000000, 80'h00000000000006000000, 80'h00000000000003000000, 80'h00000000000000800000,
    80'h00000000000000400000, 80'h00000000000000300000, 80'h00000000000000180000, 80'h000000000000000c0000,
    80'h00000000000000060000, 80'h00000000000000030000, 80'h00000000000000018000, 80'h0000000000000000c000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_138 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000018000000000, 80'h00000000008000000000, 80'h00000000004000000000, 80'h00000000002000000000,
    80'h00000000001000000000, 80'h00000000001800000000, 80'h00000000000c00000000, 80'h00000000000600000000,
    80'h00000000000300000000, 80'h00000000000180000000, 80'h000000000000c0000000, 80'h00000000000040000000,
    80'h00000000000020000000, 80'h00000000000010000000, 80'h00000000000008000000, 80'h0000000000000c000000,
    80'h00000000000006000000, 80'h00000000000003000000, 80'h00000000000001800000, 80'h00000000000000c00000,
    80'h00000000000000600000, 80'h00000000000000200000, 80'h00000000000000100000, 80'h00000000000000080000,
    80'h00000000000000040000, 80'h00000000000000060000, 80'h00000000000000030000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_144 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000008000000000, 80'h0000000000c000000000, 80'h00000000006000000000,
    80'h00000000002000000000, 80'h00000000001000000000, 80'h00000000001800000000, 80'h00000000000c00000000,
    80'h00000000000400000000, 80'h00000000000200000000, 80'h00000000000300000000, 80'h00000000000100000000,
    80'h00000000000080000000, 80'h000000000000c0000000, 80'h00000000000060000000, 80'h00000000000020000000,
    80'h00000000000010000000, 80'h00000000000018000000, 80'h0000000000000c000000, 80'h00000000000004000000,
    80'h00000000000002000000, 80'h00000000000003000000, 80'h00000000000001000000, 80'h00000000000000800000,
    80'h00000000000000c00000, 80'h00000000000000600000, 80'h00000000000000200000, 80'h00000000000000100000,
    80'h00000000000000180000, 80'h00000000000000080000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_150 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000008000000000, 80'h0000000000c000000000, 80'h00000000004000000000,
    80'h00000000006000000000, 80'h00000000002000000000, 80'h00000000003000000000, 80'h00000000001000000000,
    80'h00000000000800000000, 80'h00000000000c00000000, 80'h00000000000400000000, 80'h00000000000600000000,
    80'h00000000000200000000, 80'h00000000000100000000, 80'h00000000000100000000, 80'h00000000000080000000,
    80'h000000000000c0000000, 80'h00000000000040000000, 80'h00000000000060000000, 80'h00000000000020000000,
    80'h00000000000010000000, 80'h00000000000018000000, 80'h00000000000008000000, 80'h0000000000000c000000,
    80'h00000000000004000000, 80'h00000000000006000000, 80'h00000000000002000000, 80'h00000000000001000000,
    80'h00000000000001800000, 80'h00000000000000800000, 80'h00000000000000c00000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_156 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000008000000000, 80'h0000000000c000000000,
    80'h00000000004000000000, 80'h00000000006000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001800000000, 80'h00000000000800000000,
    80'h00000000000c00000000, 80'h00000000000400000000, 80'h00000000000600000000, 80'h00000000000200000000,
    80'h00000000000200000000, 80'h00000000000100000000, 80'h00000000000100000000, 80'h00000000000180000000,
    80'h00000000000080000000, 80'h000000000000c0000000, 80'h00000000000040000000, 80'h00000000000060000000,
    80'h00000000000020000000, 80'h00000000000020000000, 80'h00000000000010000000, 80'h00000000000010000000,
    80'h00000000000018000000, 80'h00000000000008000000, 80'h0000000000000c000000, 80'h00000000000004000000,
    80'h00000000000006000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_162 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h0000000000c000000000, 80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000006000000000,
    80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000003000000000, 80'h00000000001000000000,
    80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000000800000000, 80'h00000000000800000000,
    80'h00000000000800000000, 80'h00000000000400000000, 80'h00000000000400000000, 80'h00000000000400000000,
    80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000300000000,
    80'h00000000000100000000, 80'h00000000000100000000, 80'h00000000000180000000, 80'h00000000000080000000,
    80'h00000000000080000000, 80'h000000000000c0000000, 80'h00000000000040000000, 80'h00000000000040000000,
    80'h00000000000060000000, 80'h00000000000020000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_168 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h0000000000c000000000,
    80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000006000000000,
    80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000003000000000, 80'h00000000001000000000, 80'h00000000001000000000, 80'h00000000001000000000,
    80'h00000000001000000000, 80'h00000000001800000000, 80'h00000000000800000000, 80'h00000000000800000000,
    80'h00000000000800000000, 80'h00000000000c00000000, 80'h00000000000400000000, 80'h00000000000400000000,
    80'h00000000000400000000, 80'h00000000000400000000, 80'h00000000000600000000, 80'h00000000000200000000,
    80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000200000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_174 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000018000000000, 80'h00000000018000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h0000000000c000000000, 80'h0000000000c000000000, 80'h00000000004000000000,
    80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000004000000000,
    80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000004000000000, 80'h00000000006000000000,
    80'h00000000006000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000, 80'h00000000002000000000,
    80'h00000000003000000000, 80'h00000000003000000000, 80'h00000000001000000000, 80'h00000000001000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_180 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_186 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000030000000000, 80'h00000000030000000000, 80'h00000000020000000000, 80'h00000000020000000000,
    80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000020000000000,
    80'h00000000020000000000, 80'h00000000060000000000, 80'h00000000060000000000, 80'h00000000040000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h000000000c0000000000,
    80'h000000000c0000000000, 80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000080000000000,
    80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000080000000000,
    80'h00000000180000000000, 80'h00000000180000000000, 80'h00000000100000000000, 80'h00000000100000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_192 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000030000000000, 80'h00000000020000000000,
    80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000060000000000, 80'h00000000060000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h000000000c0000000000,
    80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000080000000000,
    80'h00000000180000000000, 80'h00000000100000000000, 80'h00000000100000000000, 80'h00000000100000000000,
    80'h00000000100000000000, 80'h00000000300000000000, 80'h00000000200000000000, 80'h00000000200000000000,
    80'h00000000200000000000, 80'h00000000600000000000, 80'h00000000400000000000, 80'h00000000400000000000,
    80'h00000000400000000000, 80'h00000000400000000000, 80'h00000000c00000000000, 80'h00000000800000000000,
    80'h00000000800000000000, 80'h00000000800000000000, 80'h00000000800000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_198 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000030000000000, 80'h00000000020000000000, 80'h00000000020000000000,
    80'h00000000060000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h000000000c0000000000,
    80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000180000000000, 80'h00000000100000000000,
    80'h00000000100000000000, 80'h00000000300000000000, 80'h00000000200000000000, 80'h00000000200000000000,
    80'h00000000600000000000, 80'h00000000400000000000, 80'h00000000400000000000, 80'h00000000400000000000,
    80'h00000000800000000000, 80'h00000000800000000000, 80'h00000000800000000000, 80'h00000001000000000000,
    80'h00000001000000000000, 80'h00000001000000000000, 80'h00000002000000000000, 80'h00000002000000000000,
    80'h00000002000000000000, 80'h00000006000000000000, 80'h00000004000000000000, 80'h00000004000000000000,
    80'h0000000c000000000000, 80'h00000008000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_204 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000060000000000,
    80'h00000000040000000000, 80'h000000000c0000000000, 80'h00000000080000000000, 80'h00000000180000000000,
    80'h00000000100000000000, 80'h00000000100000000000, 80'h00000000200000000000, 80'h00000000200000000000,
    80'h00000000600000000000, 80'h00000000400000000000, 80'h00000000c00000000000, 80'h00000000800000000000,
    80'h00000001800000000000, 80'h00000001000000000000, 80'h00000001000000000000, 80'h00000002000000000000,
    80'h00000002000000000000, 80'h00000006000000000000, 80'h00000004000000000000, 80'h0000000c000000000000,
    80'h00000008000000000000, 80'h00000018000000000000, 80'h00000010000000000000, 80'h00000010000000000000,
    80'h00000020000000000000, 80'h00000020000000000000, 80'h00000060000000000000, 80'h00000040000000000000,
    80'h00000040000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_210 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000030000000000, 80'h00000000020000000000, 80'h00000000060000000000, 80'h00000000040000000000,
    80'h000000000c0000000000, 80'h00000000080000000000, 80'h00000000100000000000, 80'h00000000300000000000,
    80'h00000000200000000000, 80'h00000000600000000000, 80'h00000000400000000000, 80'h00000000800000000000,
    80'h00000000800000000000, 80'h00000001000000000000, 80'h00000003000000000000, 80'h00000002000000000000,
    80'h00000006000000000000, 80'h00000004000000000000, 80'h00000008000000000000, 80'h00000018000000000000,
    80'h00000010000000000000, 80'h00000030000000000000, 80'h00000020000000000000, 80'h00000060000000000000,
    80'h00000040000000000000, 80'h00000080000000000000, 80'h00000180000000000000, 80'h00000100000000000000,
    80'h00000300000000000000, 80'h00000200000000000000, 80'h00000600000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_216 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000030000000000, 80'h00000000020000000000, 80'h00000000040000000000, 80'h000000000c0000000000,
    80'h00000000180000000000, 80'h00000000100000000000, 80'h00000000200000000000, 80'h00000000600000000000,
    80'h00000000c00000000000, 80'h00000000800000000000, 80'h00000001000000000000, 80'h00000003000000000000,
    80'h00000002000000000000, 80'h00000004000000000000, 80'h0000000c000000000000, 80'h00000018000000000000,
    80'h00000010000000000000, 80'h00000020000000000000, 80'h00000060000000000000, 80'h000000c0000000000000,
    80'h00000080000000000000, 80'h00000180000000000000, 80'h00000300000000000000, 80'h00000200000000000000,
    80'h00000400000000000000, 80'h00000c00000000000000, 80'h00001800000000000000, 80'h00001000000000000000,
    80'h00002000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_222 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000,
    80'h00000000030000000000, 80'h00000000060000000000, 80'h000000000c0000000000, 80'h00000000180000000000,
    80'h00000000300000000000, 80'h00000000200000000000, 80'h00000000400000000000, 80'h00000000800000000000,
    80'h00000001000000000000, 80'h00000003000000000000, 80'h00000006000000000000, 80'h0000000c000000000000,
    80'h00000018000000000000, 80'h00000030000000000000, 80'h00000060000000000000, 80'h00000040000000000000,
    80'h00000080000000000000, 80'h00000100000000000000, 80'h00000200000000000000, 80'h00000600000000000000,
    80'h00000c00000000000000, 80'h00001800000000000000, 80'h00003000000000000000, 80'h00006000000000000000,
    80'h0000c000000000000000, 80'h00008000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_228 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000,
    80'h00000000030000000000, 80'h00000000040000000000, 80'h00000000080000000000, 80'h00000000300000000000,
    80'h00000000600000000000, 80'h00000000c00000000000, 80'h00000001800000000000, 80'h00000003000000000000,
    80'h00000006000000000000, 80'h0000000c000000000000, 80'h00000010000000000000, 80'h00000020000000000000,
    80'h000000c0000000000000, 80'h00000180000000000000, 80'h00000300000000000000, 80'h00000600000000000000,
    80'h00000c00000000000000, 80'h00001800000000000000, 80'h00003000000000000000, 80'h00004000000000000000,
    80'h00008000000000000000, 80'h00030000000000000000, 80'h00060000000000000000, 80'h00040000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_234 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000,
    80'h00000000060000000000, 80'h000000000c0000000000, 80'h00000000180000000000, 80'h00000000600000000000,
    80'h00000000c00000000000, 80'h00000001800000000000, 80'h00000006000000000000, 80'h0000000c000000000000,
    80'h00000030000000000000, 80'h00000060000000000000, 80'h000000c0000000000000, 80'h00000300000000000000,
    80'h00000600000000000000, 80'h00000c00000000000000, 80'h00003000000000000000, 80'h00006000000000000000,
    80'h00018000000000000000, 80'h00030000000000000000, 80'h00060000000000000000, 80'h00180000000000000000,
    80'h00300000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_240 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000,
    80'h00000000060000000000, 80'h000000001c0000000000, 80'h00000000700000000000, 80'h00000000c00000000000,
    80'h00000003000000000000, 80'h0000000e000000000000, 80'h00000018000000000000, 80'h00000060000000000000,
    80'h00000180000000000000, 80'h00000700000000000000, 80'h00000c00000000000000, 80'h00003000000000000000,
    80'h0000e000000000000000, 80'h00038000000000000000, 80'h00060000000000000000, 80'h00180000000000000000,
    80'h00700000000000000000, 80'h00400000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_246 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000,
    80'h000000000e0000000000, 80'h00000000380000000000, 80'h00000000e00000000000, 80'h00000007000000000000,
    80'h0000001c000000000000, 80'h00000070000000000000, 80'h000001c0000000000000, 80'h00000e00000000000000,
    80'h00003800000000000000, 80'h0000e000000000000000, 80'h00038000000000000000, 80'h001c0000000000000000,
    80'h00700000000000000000, 80'h01c00000000000000000, 80'h01000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_252 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000,
    80'h000000001e0000000000, 80'h00000000f00000000000, 80'h00000007800000000000, 80'h0000003c000000000000,
    80'h000001c0000000000000, 80'h00000e00000000000000, 80'h0000f000000000000000, 80'h00078000000000000000,
    80'h003c0000000000000000, 80'h01e00000000000000000, 80'h03000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_258 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000078000000000,
    80'h00000000fc0000000000, 80'h0000000f800000000000, 80'h000001f8000000000000, 80'h00003f00000000000000,
    80'h0003e000000000000000, 80'h007e0000000000000000, 80'h07c00000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_264 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h000000003f8000000000,
    80'h0000007ff00000000000, 80'h0001ffe0000000000000, 80'h03ff8000000000000000, 80'h0f000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_270 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0fffffffff8000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_276 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0f000000000000000000,
    80'h03ff8000000000000000, 80'h0001ffe0000000000000, 80'h0000007ff00000000000, 80'h000000003f8000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_282 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h07c00000000000000000, 80'h007e0000000000000000, 80'h0003e000000000000000, 80'h00003f00000000000000,
    80'h000001f8000000000000, 80'h0000000fc00000000000, 80'h00000000fc0000000000, 80'h00000000078000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_288 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h03000000000000000000, 80'h01e00000000000000000, 80'h003c0000000000000000, 80'h00038000000000000000,
    80'h00007000000000000000, 80'h00000f00000000000000, 80'h000001e0000000000000, 80'h0000003c000000000000,
    80'h00000007800000000000, 80'h00000000f00000000000, 80'h000000001e0000000000, 80'h00000000038000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_294 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h01c00000000000000000, 80'h00700000000000000000, 80'h000e0000000000000000,
    80'h00038000000000000000, 80'h0000e000000000000000, 80'h00003800000000000000, 80'h00000700000000000000,
    80'h000001c0000000000000, 80'h00000070000000000000, 80'h0000001c000000000000, 80'h00000003800000000000,
    80'h00000000e00000000000, 80'h00000000380000000000, 80'h000000000e0000000000, 80'h00000000018000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_300 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00400000000000000000, 80'h00700000000000000000, 80'h001c0000000000000000,
    80'h00060000000000000000, 80'h00018000000000000000, 80'h0000e000000000000000, 80'h00003800000000000000,
    80'h00000c00000000000000, 80'h00000300000000000000, 80'h000001c0000000000000, 80'h00000060000000000000,
    80'h00000018000000000000, 80'h00000006000000000000, 80'h00000003800000000000, 80'h00000000c00000000000,
    80'h00000000300000000000, 80'h000000001c0000000000, 80'h00000000070000000000, 80'h00000000018000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_306 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00100000000000000000, 80'h000c0000000000000000,
    80'h00060000000000000000, 80'h00030000000000000000, 80'h0000c000000000000000, 80'h00006000000000000000,
    80'h00003800000000000000, 80'h00000c00000000000000, 80'h00000600000000000000, 80'h00000180000000000000,
    80'h000000c0000000000000, 80'h00000060000000000000, 80'h00000018000000000000, 80'h0000000c000000000000,
    80'h00000003000000000000, 80'h00000001800000000000, 80'h00000000c00000000000, 80'h00000000300000000000,
    80'h00000000180000000000, 80'h000000000c0000000000, 80'h00000000030000000000, 80'h00000000018000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_312 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00030000000000000000, 80'h00018000000000000000, 80'h0000c000000000000000, 80'h00006000000000000000,
    80'h00003000000000000000, 80'h00001800000000000000, 80'h00000c00000000000000, 80'h00000200000000000000,
    80'h00000100000000000000, 80'h000000c0000000000000, 80'h00000060000000000000, 80'h00000030000000000000,
    80'h00000018000000000000, 80'h0000000c000000000000, 80'h00000006000000000000, 80'h00000003000000000000,
    80'h00000000800000000000, 80'h00000000400000000000, 80'h00000000300000000000, 80'h00000000180000000000,
    80'h000000000c0000000000, 80'h00000000060000000000, 80'h00000000030000000000, 80'h00000000018000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_318 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h0000c000000000000000, 80'h00006000000000000000, 80'h00002000000000000000,
    80'h00001000000000000000, 80'h00000800000000000000, 80'h00000400000000000000, 80'h00000600000000000000,
    80'h00000300000000000000, 80'h00000180000000000000, 80'h000000c0000000000000, 80'h00000060000000000000,
    80'h00000030000000000000, 80'h00000010000000000000, 80'h00000008000000000000, 80'h00000004000000000000,
    80'h00000002000000000000, 80'h00000003000000000000, 80'h00000001800000000000, 80'h00000000c00000000000,
    80'h00000000600000000000, 80'h00000000300000000000, 80'h00000000180000000000, 80'h00000000080000000000,
    80'h00000000040000000000, 80'h00000000020000000000, 80'h00000000010000000000, 80'h00000000018000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_324 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00001000000000000000, 80'h00001800000000000000,
    80'h00000800000000000000, 80'h00000400000000000000, 80'h00000600000000000000, 80'h00000300000000000000,
    80'h00000100000000000000, 80'h00000080000000000000, 80'h000000c0000000000000, 80'h00000040000000000000,
    80'h00000020000000000000, 80'h00000030000000000000, 80'h00000018000000000000, 80'h00000008000000000000,
    80'h00000004000000000000, 80'h00000006000000000000, 80'h00000003000000000000, 80'h00000001000000000000,
    80'h00000000800000000000, 80'h00000000c00000000000, 80'h00000000400000000000, 80'h00000000200000000000,
    80'h00000000300000000000, 80'h00000000180000000000, 80'h00000000080000000000, 80'h00000000040000000000,
    80'h00000000060000000000, 80'h00000000030000000000, 80'h00000000010000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_330 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000300000000000000, 80'h00000100000000000000, 80'h00000180000000000000,
    80'h00000080000000000000, 80'h00000040000000000000, 80'h00000060000000000000, 80'h00000020000000000000,
    80'h00000030000000000000, 80'h00000010000000000000, 80'h00000018000000000000, 80'h00000008000000000000,
    80'h00000004000000000000, 80'h00000006000000000000, 80'h00000002000000000000, 80'h00000003000000000000,
    80'h00000001000000000000, 80'h00000000800000000000, 80'h00000000800000000000, 80'h00000000400000000000,
    80'h00000000600000000000, 80'h00000000200000000000, 80'h00000000300000000000, 80'h00000000100000000000,
    80'h00000000080000000000, 80'h000000000c0000000000, 80'h00000000040000000000, 80'h00000000060000000000,
    80'h00000000020000000000, 80'h00000000030000000000, 80'h00000000010000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_336 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000060000000000000,
    80'h00000020000000000000, 80'h00000030000000000000, 80'h00000010000000000000, 80'h00000018000000000000,
    80'h00000008000000000000, 80'h00000008000000000000, 80'h00000004000000000000, 80'h00000004000000000000,
    80'h00000006000000000000, 80'h00000002000000000000, 80'h00000003000000000000, 80'h00000001000000000000,
    80'h00000001800000000000, 80'h00000000800000000000, 80'h00000000800000000000, 80'h00000000400000000000,
    80'h00000000400000000000, 80'h00000000600000000000, 80'h00000000200000000000, 80'h00000000300000000000,
    80'h00000000100000000000, 80'h00000000180000000000, 80'h00000000080000000000, 80'h00000000080000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000060000000000, 80'h00000000020000000000,
    80'h00000000030000000000, 80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_342 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000004000000000000, 80'h00000006000000000000,
    80'h00000002000000000000, 80'h00000002000000000000, 80'h00000003000000000000, 80'h00000001000000000000,
    80'h00000001000000000000, 80'h00000001800000000000, 80'h00000000800000000000, 80'h00000000800000000000,
    80'h00000000c00000000000, 80'h00000000400000000000, 80'h00000000400000000000, 80'h00000000400000000000,
    80'h00000000200000000000, 80'h00000000200000000000, 80'h00000000200000000000, 80'h00000000100000000000,
    80'h00000000100000000000, 80'h00000000100000000000, 80'h00000000080000000000, 80'h00000000080000000000,
    80'h00000000080000000000, 80'h000000000c0000000000, 80'h00000000040000000000, 80'h00000000040000000000,
    80'h00000000060000000000, 80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000030000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_348 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000400000000000, 80'h00000000400000000000, 80'h00000000400000000000,
    80'h00000000400000000000, 80'h00000000600000000000, 80'h00000000200000000000, 80'h00000000200000000000,
    80'h00000000200000000000, 80'h00000000200000000000, 80'h00000000300000000000, 80'h00000000100000000000,
    80'h00000000100000000000, 80'h00000000100000000000, 80'h00000000180000000000, 80'h00000000080000000000,
    80'h00000000080000000000, 80'h00000000080000000000, 80'h00000000080000000000, 80'h000000000c0000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000,
    80'h00000000060000000000, 80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000020000000000,
    80'h00000000030000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] second_354 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000080000000000, 80'h00000000080000000000, 80'h000000000c0000000000, 80'h000000000c0000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000,
    80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000040000000000, 80'h00000000060000000000,
    80'h00000000060000000000, 80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000020000000000,
    80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000020000000000, 80'h00000000020000000000,
    80'h00000000020000000000, 80'h00000000030000000000, 80'h00000000030000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000010000000000,
    80'h00000000010000000000, 80'h00000000010000000000, 80'h00000000018000000000, 80'h00000000018000000000,
    80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000, 80'h00000000008000000000,
    80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};


wire [0:79] minute_000 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_006 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000003800000000, 80'h00000000003800000000, 80'h00000000003800000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_012 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000400000000, 80'h00000000000e00000000, 80'h00000000000e00000000,
    80'h00000000000e00000000, 80'h00000000000e00000000, 80'h00000000000e00000000, 80'h00000000001c00000000,
    80'h00000000001c00000000, 80'h00000000001c00000000, 80'h00000000001c00000000, 80'h00000000003c00000000,
    80'h00000000003800000000, 80'h00000000003800000000, 80'h00000000003800000000, 80'h00000000003800000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000,
    80'h00000000007000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_018 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000180000000, 80'h000000000001c0000000,
    80'h000000000001c0000000, 80'h00000000000380000000, 80'h00000000000380000000, 80'h00000000000380000000,
    80'h00000000000700000000, 80'h00000000000700000000, 80'h00000000000700000000, 80'h00000000000e00000000,
    80'h00000000000e00000000, 80'h00000000000e00000000, 80'h00000000001c00000000, 80'h00000000001c00000000,
    80'h00000000001c00000000, 80'h00000000003c00000000, 80'h00000000003800000000, 80'h00000000003800000000,
    80'h00000000007800000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h0000000000f000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000001e000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_024 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000020000000,
    80'h00000000000078000000, 80'h00000000000070000000, 80'h000000000000f0000000, 80'h000000000000e0000000,
    80'h000000000000e0000000, 80'h000000000001c0000000, 80'h000000000001c0000000, 80'h000000000003c0000000,
    80'h00000000000380000000, 80'h00000000000780000000, 80'h00000000000700000000, 80'h00000000000f00000000,
    80'h00000000000e00000000, 80'h00000000000e00000000, 80'h00000000001c00000000, 80'h00000000001c00000000,
    80'h00000000003c00000000, 80'h00000000003800000000, 80'h00000000007800000000, 80'h00000000007000000000,
    80'h0000000000f000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_030 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000008000000, 80'h0000000000000e000000, 80'h0000000000001e000000, 80'h0000000000001c000000,
    80'h0000000000003c000000, 80'h00000000000038000000, 80'h00000000000070000000, 80'h000000000000f0000000,
    80'h000000000000e0000000, 80'h000000000001e0000000, 80'h000000000001c0000000, 80'h000000000003c0000000,
    80'h00000000000780000000, 80'h00000000000700000000, 80'h00000000000f00000000, 80'h00000000000e00000000,
    80'h00000000001e00000000, 80'h00000000001c00000000, 80'h00000000003800000000, 80'h00000000007800000000,
    80'h00000000007000000000, 80'h0000000000f000000000, 80'h0000000000e000000000, 80'h0000000001e000000000,
    80'h0000000003c000000000, 80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_036 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000003000000, 80'h00000000000003800000,
    80'h00000000000007800000, 80'h0000000000000f000000, 80'h0000000000001e000000, 80'h0000000000001c000000,
    80'h0000000000003c000000, 80'h00000000000078000000, 80'h00000000000070000000, 80'h000000000000f0000000,
    80'h000000000001e0000000, 80'h000000000003c0000000, 80'h00000000000380000000, 80'h00000000000780000000,
    80'h00000000000f00000000, 80'h00000000001e00000000, 80'h00000000001c00000000, 80'h00000000003c00000000,
    80'h00000000007800000000, 80'h00000000007000000000, 80'h0000000000f000000000, 80'h0000000001e000000000,
    80'h0000000003c000000000, 80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_042 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000e00000, 80'h00000000000001e00000, 80'h00000000000003c00000, 80'h00000000000003c00000,
    80'h00000000000007800000, 80'h0000000000000f000000, 80'h0000000000001e000000, 80'h0000000000003c000000,
    80'h00000000000078000000, 80'h000000000000f0000000, 80'h000000000001e0000000, 80'h000000000003c0000000,
    80'h00000000000780000000, 80'h00000000000780000000, 80'h00000000000f00000000, 80'h00000000001e00000000,
    80'h00000000003c00000000, 80'h00000000007800000000, 80'h0000000000f000000000, 80'h0000000001e000000000,
    80'h0000000003c000000000, 80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_048 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000100000, 80'h00000000000000380000, 80'h00000000000000780000,
    80'h00000000000000f00000, 80'h00000000000001e00000, 80'h00000000000007c00000, 80'h0000000000000f800000,
    80'h0000000000001f000000, 80'h0000000000003e000000, 80'h0000000000007c000000, 80'h000000000000f0000000,
    80'h000000000001e0000000, 80'h000000000003c0000000, 80'h00000000000780000000, 80'h00000000000f00000000,
    80'h00000000003e00000000, 80'h00000000007c00000000, 80'h0000000000f800000000, 80'h0000000001f000000000,
    80'h0000000003c000000000, 80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_054 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h000000000000000c0000, 80'h000000000000003e0000, 80'h000000000000007c0000, 80'h00000000000000f80000,
    80'h00000000000003e00000, 80'h00000000000007c00000, 80'h0000000000001f000000, 80'h0000000000003e000000,
    80'h0000000000007c000000, 80'h000000000001f0000000, 80'h000000000003e0000000, 80'h00000000000fc0000000,
    80'h00000000001f00000000, 80'h00000000003e00000000, 80'h0000000000f800000000, 80'h0000000001f000000000,
    80'h0000000003e000000000, 80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_060 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000060000, 80'h000000000000000f0000,
    80'h000000000000003f0000, 80'h00000000000000fc0000, 80'h00000000000003f00000, 80'h00000000000007e00000,
    80'h0000000000001f800000, 80'h0000000000007e000000, 80'h000000000000fc000000, 80'h000000000003f0000000,
    80'h00000000000fc0000000, 80'h00000000003f00000000, 80'h00000000007e00000000, 80'h0000000001f800000000,
    80'h0000000003e000000000, 80'h00000000018000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_066 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000010000, 80'h00000000000000078000, 80'h000000000000001f8000, 80'h000000000000007f0000,
    80'h00000000000003fc0000, 80'h0000000000000ff00000, 80'h0000000000003f800000, 80'h000000000000fe000000,
    80'h000000000007f8000000, 80'h00000000001fe0000000, 80'h00000000007f00000000, 80'h0000000001fc00000000,
    80'h0000000003f000000000, 80'h0000000003c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_072 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000000000001c000,
    80'h000000000000000fc000, 80'h000000000000007fc000, 80'h00000000000003fe0000, 80'h0000000000001ff00000,
    80'h000000000000ff800000, 80'h00000000000ffc000000, 80'h00000000007fe0000000, 80'h0000000003ff00000000,
    80'h0000000003f800000000, 80'h0000000003c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_078 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000004000, 80'h0000000000000007c000, 80'h00000000000000ffe000,
    80'h0000000000000fffc000, 80'h000000000001fff80000, 80'h00000000003fff800000, 80'h0000000003fff0000000,
    80'h0000000003fe00000000, 80'h0000000003e000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_084 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h0000000000000000e000, 80'h00000000000003ffe000, 80'h000000000007ffffe000, 80'h0000000003ffffff0000,
    80'h0000000003fffc000000, 80'h0000000003f800000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_090 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003ffffffe000,
    80'h0000000003ffffffe000, 80'h0000000003ffffffe000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_096 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003f800000000,
    80'h0000000003fffc000000, 80'h0000000003ffffff0000, 80'h000000000007ffffe000, 80'h00000000000003ffe000,
    80'h0000000000000000e000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_102 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003c000000000,
    80'h0000000003fe00000000, 80'h0000000003fff0000000, 80'h00000000003fff800000, 80'h000000000001fff80000,
    80'h0000000000000fffc000, 80'h00000000000000ffe000, 80'h0000000000000007c000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_108 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003c000000000,
    80'h0000000003f800000000, 80'h0000000003ff00000000, 80'h00000000007fe0000000, 80'h00000000000ffc000000,
    80'h000000000001ff800000, 80'h0000000000003ff00000, 80'h00000000000003fe0000, 80'h000000000000007fc000,
    80'h000000000000000fc000, 80'h00000000000000018000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_114 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000,
    80'h0000000003f000000000, 80'h0000000003fc00000000, 80'h00000000007f00000000, 80'h00000000001fc0000000,
    80'h000000000007f8000000, 80'h000000000001fe000000, 80'h0000000000003f800000, 80'h0000000000000fe00000,
    80'h00000000000003fc0000, 80'h00000000000000ff0000, 80'h000000000000001f8000, 80'h00000000000000070000,
    80'h00000000000000010000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_120 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000, 80'h00000000038000000000,
    80'h0000000003e000000000, 80'h0000000001f800000000, 80'h0000000000fc00000000, 80'h00000000003f00000000,
    80'h00000000000fc0000000, 80'h000000000003f0000000, 80'h000000000001f8000000, 80'h0000000000007e000000,
    80'h0000000000001f800000, 80'h0000000000000fc00000, 80'h00000000000003f00000, 80'h00000000000000fc0000,
    80'h000000000000003f0000, 80'h000000000000001e0000, 80'h00000000000000060000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_126 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000, 80'h00000000038000000000,
    80'h0000000003c000000000, 80'h0000000001f000000000, 80'h0000000000f800000000, 80'h00000000007e00000000,
    80'h00000000001f00000000, 80'h00000000000f80000000, 80'h000000000003e0000000, 80'h000000000001f0000000,
    80'h000000000000f8000000, 80'h0000000000003e000000, 80'h0000000000001f000000, 80'h0000000000000fc00000,
    80'h00000000000003e00000, 80'h00000000000001f00000, 80'h000000000000007c0000, 80'h000000000000003c0000,
    80'h00000000000000180000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_132 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000, 80'h00000000038000000000,
    80'h0000000003c000000000, 80'h0000000001e000000000, 80'h0000000000f000000000, 80'h00000000007800000000,
    80'h00000000003c00000000, 80'h00000000001f00000000, 80'h00000000000f80000000, 80'h000000000007c0000000,
    80'h000000000003e0000000, 80'h000000000000f0000000, 80'h00000000000078000000, 80'h0000000000003c000000,
    80'h0000000000001e000000, 80'h0000000000000f000000, 80'h00000000000007c00000, 80'h00000000000003e00000,
    80'h00000000000001f00000, 80'h00000000000000f00000, 80'h00000000000000300000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_138 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000, 80'h00000000038000000000,
    80'h0000000003c000000000, 80'h0000000001e000000000, 80'h0000000000f000000000, 80'h0000000000f000000000,
    80'h00000000007800000000, 80'h00000000003c00000000, 80'h00000000001e00000000, 80'h00000000000f00000000,
    80'h00000000000780000000, 80'h000000000003c0000000, 80'h000000000001e0000000, 80'h000000000000f0000000,
    80'h00000000000078000000, 80'h0000000000007c000000, 80'h0000000000003c000000, 80'h0000000000001e000000,
    80'h0000000000000f000000, 80'h00000000000007800000, 80'h00000000000003c00000, 80'h00000000000001e00000,
    80'h00000000000000c00000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_144 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000, 80'h00000000038000000000,
    80'h0000000003c000000000, 80'h0000000001c000000000, 80'h0000000001e000000000, 80'h0000000000f000000000,
    80'h00000000007800000000, 80'h00000000003800000000, 80'h00000000003c00000000, 80'h00000000001e00000000,
    80'h00000000000e00000000, 80'h00000000000f00000000, 80'h00000000000780000000, 80'h000000000003c0000000,
    80'h000000000001c0000000, 80'h000000000001e0000000, 80'h000000000000f0000000, 80'h00000000000070000000,
    80'h00000000000038000000, 80'h0000000000003c000000, 80'h0000000000001e000000, 80'h0000000000000e000000,
    80'h0000000000000f000000, 80'h00000000000007000000, 80'h00000000000002000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_150 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000010000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h0000000001c000000000, 80'h0000000001e000000000, 80'h0000000000e000000000,
    80'h0000000000f000000000, 80'h00000000007000000000, 80'h00000000007800000000, 80'h00000000003800000000,
    80'h00000000001c00000000, 80'h00000000001e00000000, 80'h00000000000e00000000, 80'h00000000000f00000000,
    80'h00000000000700000000, 80'h00000000000780000000, 80'h000000000003c0000000, 80'h000000000001c0000000,
    80'h000000000001e0000000, 80'h000000000000e0000000, 80'h000000000000f0000000, 80'h00000000000070000000,
    80'h00000000000038000000, 80'h0000000000003c000000, 80'h0000000000001c000000, 80'h00000000000018000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_156 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000030000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h0000000003c000000000, 80'h0000000001c000000000, 80'h0000000001e000000000,
    80'h0000000000e000000000, 80'h0000000000f000000000, 80'h00000000007000000000, 80'h00000000007000000000,
    80'h00000000003800000000, 80'h00000000003800000000, 80'h00000000003c00000000, 80'h00000000001c00000000,
    80'h00000000001e00000000, 80'h00000000000e00000000, 80'h00000000000f00000000, 80'h00000000000700000000,
    80'h00000000000700000000, 80'h00000000000380000000, 80'h00000000000380000000, 80'h000000000003c0000000,
    80'h000000000001c0000000, 80'h000000000001e0000000, 80'h000000000000e0000000, 80'h000000000000f0000000,
    80'h00000000000060000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_162 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h0000000003c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000003800000000,
    80'h00000000003800000000, 80'h00000000003800000000, 80'h00000000001c00000000, 80'h00000000001c00000000,
    80'h00000000001c00000000, 80'h00000000000e00000000, 80'h00000000000e00000000, 80'h00000000000e00000000,
    80'h00000000000700000000, 80'h00000000000700000000, 80'h00000000000700000000, 80'h00000000000380000000,
    80'h00000000000380000000, 80'h00000000000380000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_168 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h0000000003c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000000e000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000,
    80'h00000000007800000000, 80'h00000000003800000000, 80'h00000000003800000000, 80'h00000000003800000000,
    80'h00000000003800000000, 80'h00000000001c00000000, 80'h00000000001c00000000, 80'h00000000001c00000000,
    80'h00000000001c00000000, 80'h00000000001e00000000, 80'h00000000000800000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_174 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000, 80'h0000000000e000000000,
    80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000007000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_180 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_186 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h000000001c0000000000, 80'h000000001c0000000000, 80'h000000001c0000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_192 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h000000000e0000000000,
    80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h000000001c0000000000, 80'h000000001c0000000000, 80'h000000001c0000000000, 80'h000000001c0000000000,
    80'h000000003c0000000000, 80'h00000000380000000000, 80'h00000000380000000000, 80'h00000000380000000000,
    80'h00000000380000000000, 80'h00000000700000000000, 80'h00000000700000000000, 80'h00000000700000000000,
    80'h00000000700000000000, 80'h00000000700000000000, 80'h00000000200000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_198 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000078000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h000000000f0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000001e0000000000,
    80'h000000001c0000000000, 80'h000000001c0000000000, 80'h000000003c0000000000, 80'h00000000380000000000,
    80'h00000000380000000000, 80'h00000000380000000000, 80'h00000000700000000000, 80'h00000000700000000000,
    80'h00000000700000000000, 80'h00000000e00000000000, 80'h00000000e00000000000, 80'h00000000e00000000000,
    80'h00000001c00000000000, 80'h00000001c00000000000, 80'h00000001c00000000000, 80'h00000003800000000000,
    80'h00000003800000000000, 80'h00000001800000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_204 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h000000000f0000000000,
    80'h000000000e0000000000, 80'h000000001e0000000000, 80'h000000001c0000000000, 80'h000000003c0000000000,
    80'h00000000380000000000, 80'h00000000380000000000, 80'h00000000700000000000, 80'h00000000700000000000,
    80'h00000000f00000000000, 80'h00000000e00000000000, 80'h00000001e00000000000, 80'h00000001c00000000000,
    80'h00000003c00000000000, 80'h00000003800000000000, 80'h00000003800000000000, 80'h00000007000000000000,
    80'h00000007000000000000, 80'h0000000f000000000000, 80'h0000000e000000000000, 80'h0000001e000000000000,
    80'h00000004000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_210 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000, 80'h0000000003c000000000,
    80'h00000000078000000000, 80'h00000000070000000000, 80'h000000000f0000000000, 80'h000000000e0000000000,
    80'h000000001e0000000000, 80'h000000001c0000000000, 80'h00000000380000000000, 80'h00000000780000000000,
    80'h00000000700000000000, 80'h00000000f00000000000, 80'h00000000e00000000000, 80'h00000001e00000000000,
    80'h00000003c00000000000, 80'h00000003800000000000, 80'h00000007800000000000, 80'h00000007000000000000,
    80'h0000000f000000000000, 80'h0000000e000000000000, 80'h0000001c000000000000, 80'h0000003c000000000000,
    80'h00000038000000000000, 80'h00000078000000000000, 80'h00000070000000000000, 80'h00000010000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_216 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000, 80'h0000000003c000000000,
    80'h00000000078000000000, 80'h000000000f0000000000, 80'h000000000e0000000000, 80'h000000001e0000000000,
    80'h000000003c0000000000, 80'h00000000380000000000, 80'h00000000780000000000, 80'h00000000f00000000000,
    80'h00000001e00000000000, 80'h00000001c00000000000, 80'h00000003c00000000000, 80'h00000007800000000000,
    80'h0000000f000000000000, 80'h0000000e000000000000, 80'h0000001e000000000000, 80'h0000003c000000000000,
    80'h00000038000000000000, 80'h00000078000000000000, 80'h000000f0000000000000, 80'h000001e0000000000000,
    80'h000001c0000000000000, 80'h000000c0000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_222 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000, 80'h0000000003c000000000,
    80'h00000000078000000000, 80'h000000000f0000000000, 80'h000000001e0000000000, 80'h000000003c0000000000,
    80'h00000000780000000000, 80'h00000000f00000000000, 80'h00000001e00000000000, 80'h00000001e00000000000,
    80'h00000003c00000000000, 80'h00000007800000000000, 80'h0000000f000000000000, 80'h0000001e000000000000,
    80'h0000003c000000000000, 80'h00000078000000000000, 80'h000000f0000000000000, 80'h000001e0000000000000,
    80'h000003c0000000000000, 80'h000003c0000000000000, 80'h00000780000000000000, 80'h00000700000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_228 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000, 80'h0000000003c000000000,
    80'h000000000f8000000000, 80'h000000001f0000000000, 80'h000000003e0000000000, 80'h000000007c0000000000,
    80'h00000000f00000000000, 80'h00000001e00000000000, 80'h00000003c00000000000, 80'h00000007800000000000,
    80'h0000000f000000000000, 80'h0000003e000000000000, 80'h0000007c000000000000, 80'h000000f8000000000000,
    80'h000001f0000000000000, 80'h000003e0000000000000, 80'h00000780000000000000, 80'h00000f00000000000000,
    80'h00001e00000000000000, 80'h00001c00000000000000, 80'h00000800000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_234 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000, 80'h0000000007c000000000,
    80'h000000000f8000000000, 80'h000000001f0000000000, 80'h000000007c0000000000, 80'h00000000f80000000000,
    80'h00000003f00000000000, 80'h00000007c00000000000, 80'h0000000f800000000000, 80'h0000003e000000000000,
    80'h0000007c000000000000, 80'h000000f8000000000000, 80'h000003e0000000000000, 80'h000007c0000000000000,
    80'h00001f00000000000000, 80'h00003e00000000000000, 80'h00007c00000000000000, 80'h00003000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_240 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000018000000000, 80'h0000000007c000000000,
    80'h000000001f8000000000, 80'h000000007e0000000000, 80'h00000000fc0000000000, 80'h00000003f00000000000,
    80'h0000000fc00000000000, 80'h0000003f000000000000, 80'h0000007e000000000000, 80'h000001f8000000000000,
    80'h000007e0000000000000, 80'h00000fc0000000000000, 80'h00003f00000000000000, 80'h0000fc00000000000000,
    80'h0000f000000000000000, 80'h00006000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_246 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003c000000000, 80'h000000000fc000000000,
    80'h000000003f8000000000, 80'h00000000fe0000000000, 80'h00000007f80000000000, 80'h0000001fe00000000000,
    80'h0000007f000000000000, 80'h000001fc000000000000, 80'h00000ff0000000000000, 80'h00003fc0000000000000,
    80'h0000fe00000000000000, 80'h0001f800000000000000, 80'h0001e000000000000000, 80'h00008000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_252 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000003c000000000, 80'h000000001fc000000000,
    80'h00000000ffc000000000, 80'h00000007fe0000000000, 80'h0000003ff00000000000, 80'h000001ff000000000000,
    80'h00000ff8000000000000, 80'h00007fc0000000000000, 80'h0003fe00000000000000, 80'h0003f000000000000000,
    80'h00038000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_258 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h0000000007c000000000, 80'h000000007fc000000000,
    80'h0000000fffc000000000, 80'h000001fffc0000000000, 80'h00001fff800000000000, 80'h0003fff0000000000000,
    80'h0007ff00000000000000, 80'h0003e000000000000000, 80'h00020000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_264 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h000000001fc000000000, 80'h0000003fffc000000000,
    80'h0000ffffffc000000000, 80'h0007ffffe00000000000, 80'h0007ffc0000000000000, 80'h00070000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_270 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h0007ffffffc000000000, 80'h0007ffffffc000000000,
    80'h0007ffffffc000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_276 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00070000000000000000,
    80'h0007ffc0000000000000, 80'h0007ffffe00000000000, 80'h0000ffffffc000000000, 80'h0000003fffc000000000,
    80'h000000001fc000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_282 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h0003e000000000000000, 80'h0007ff00000000000000, 80'h0003fff0000000000000,
    80'h00001fff800000000000, 80'h000001fffc0000000000, 80'h0000000fffc000000000, 80'h000000007fc000000000,
    80'h0000000003c000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_288 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00018000000000000000, 80'h0003f000000000000000,
    80'h0003fe00000000000000, 80'h00007fc0000000000000, 80'h00000ffc000000000000, 80'h000001ff800000000000,
    80'h0000003ff00000000000, 80'h00000007fe0000000000, 80'h00000000ffc000000000, 80'h000000001fc000000000,
    80'h0000000003c000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_294 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00008000000000000000,
    80'h0000e000000000000000, 80'h0001f800000000000000, 80'h0000ff00000000000000, 80'h00003fc0000000000000,
    80'h000007f0000000000000, 80'h000001fc000000000000, 80'h0000007f800000000000, 80'h0000001fe00000000000,
    80'h00000003f80000000000, 80'h00000000fe0000000000, 80'h000000003fc000000000, 80'h000000000fc000000000,
    80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_300 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00006000000000000000, 80'h00007800000000000000, 80'h0000fc00000000000000,
    80'h00003f00000000000000, 80'h00000fc0000000000000, 80'h000003f0000000000000, 80'h000001f8000000000000,
    80'h0000007e000000000000, 80'h0000001f800000000000, 80'h0000000fc00000000000, 80'h00000003f00000000000,
    80'h00000000fc0000000000, 80'h000000003f0000000000, 80'h000000001f8000000000, 80'h0000000007c000000000,
    80'h0000000001c000000000, 80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_306 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00001800000000000000,
    80'h00003c00000000000000, 80'h00003e00000000000000, 80'h00000f80000000000000, 80'h000007c0000000000000,
    80'h000003f0000000000000, 80'h000000f8000000000000, 80'h0000007c000000000000, 80'h0000001f000000000000,
    80'h0000000f800000000000, 80'h00000007c00000000000, 80'h00000001f00000000000, 80'h00000000f80000000000,
    80'h000000007e0000000000, 80'h000000001f0000000000, 80'h000000000f8000000000, 80'h0000000003c000000000,
    80'h0000000001c000000000, 80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_312 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000c00000000000000, 80'h00000f00000000000000, 80'h00000f80000000000000,
    80'h000007c0000000000000, 80'h000003e0000000000000, 80'h000000f0000000000000, 80'h00000078000000000000,
    80'h0000003c000000000000, 80'h0000001e000000000000, 80'h0000000f000000000000, 80'h00000007c00000000000,
    80'h00000003e00000000000, 80'h00000001f00000000000, 80'h00000000f80000000000, 80'h000000003c0000000000,
    80'h000000001e0000000000, 80'h000000000f0000000000, 80'h00000000078000000000, 80'h0000000003c000000000,
    80'h0000000001c000000000, 80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_318 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000300000000000000,
    80'h00000780000000000000, 80'h000003c0000000000000, 80'h000001e0000000000000, 80'h000000f0000000000000,
    80'h00000078000000000000, 80'h0000003c000000000000, 80'h0000003e000000000000, 80'h0000001e000000000000,
    80'h0000000f000000000000, 80'h00000007800000000000, 80'h00000003c00000000000, 80'h00000001e00000000000,
    80'h00000000f00000000000, 80'h00000000780000000000, 80'h000000003c0000000000, 80'h000000001e0000000000,
    80'h000000000f0000000000, 80'h000000000f0000000000, 80'h00000000078000000000, 80'h0000000003c000000000,
    80'h0000000001c000000000, 80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_324 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000040000000000000, 80'h000000e0000000000000, 80'h000000f0000000000000,
    80'h00000070000000000000, 80'h00000078000000000000, 80'h0000003c000000000000, 80'h0000001c000000000000,
    80'h0000000e000000000000, 80'h0000000f000000000000, 80'h00000007800000000000, 80'h00000003800000000000,
    80'h00000003c00000000000, 80'h00000001e00000000000, 80'h00000000f00000000000, 80'h00000000700000000000,
    80'h00000000780000000000, 80'h000000003c0000000000, 80'h000000001c0000000000, 80'h000000001e0000000000,
    80'h000000000f0000000000, 80'h00000000078000000000, 80'h00000000038000000000, 80'h0000000003c000000000,
    80'h0000000001c000000000, 80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_330 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000018000000000000, 80'h00000038000000000000, 80'h0000003c000000000000, 80'h0000001c000000000000,
    80'h0000000e000000000000, 80'h0000000f000000000000, 80'h00000007000000000000, 80'h00000007800000000000,
    80'h00000003800000000000, 80'h00000003c00000000000, 80'h00000001e00000000000, 80'h00000000e00000000000,
    80'h00000000f00000000000, 80'h00000000700000000000, 80'h00000000780000000000, 80'h00000000380000000000,
    80'h000000001c0000000000, 80'h000000001e0000000000, 80'h000000000e0000000000, 80'h000000000f0000000000,
    80'h00000000070000000000, 80'h00000000078000000000, 80'h00000000038000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h00000000008000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_336 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000006000000000000,
    80'h0000000f000000000000, 80'h00000007000000000000, 80'h00000007800000000000, 80'h00000003800000000000,
    80'h00000003c00000000000, 80'h00000001c00000000000, 80'h00000001c00000000000, 80'h00000000e00000000000,
    80'h00000000e00000000000, 80'h00000000f00000000000, 80'h00000000700000000000, 80'h00000000780000000000,
    80'h00000000380000000000, 80'h000000003c0000000000, 80'h000000001c0000000000, 80'h000000001c0000000000,
    80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000f0000000000, 80'h00000000070000000000,
    80'h00000000078000000000, 80'h00000000038000000000, 80'h0000000003c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000000c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_342 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000001c00000000000, 80'h00000001c00000000000,
    80'h00000001c00000000000, 80'h00000000e00000000000, 80'h00000000e00000000000, 80'h00000000e00000000000,
    80'h00000000700000000000, 80'h00000000700000000000, 80'h00000000700000000000, 80'h00000000380000000000,
    80'h00000000380000000000, 80'h00000000380000000000, 80'h000000001c0000000000, 80'h000000001c0000000000,
    80'h000000001c0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000078000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h0000000003c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_348 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000100000000000, 80'h00000000780000000000, 80'h00000000380000000000,
    80'h00000000380000000000, 80'h00000000380000000000, 80'h00000000380000000000, 80'h000000001c0000000000,
    80'h000000001c0000000000, 80'h000000001c0000000000, 80'h000000001c0000000000, 80'h000000001e0000000000,
    80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h00000000070000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h0000000003c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};

wire [0:79] minute_354 [0:79] = '{
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h000000000e0000000000, 80'h000000000e0000000000, 80'h000000000e0000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000070000000000,
    80'h00000000070000000000, 80'h00000000070000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000,
    80'h00000000038000000000, 80'h00000000038000000000, 80'h00000000038000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000, 80'h0000000001c000000000,
    80'h0000000001c000000000, 80'h0000000001c000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000,
    80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000, 80'h00000000000000000000
};


wire [0:79] clock [0:79] = '{
    80'h00000003ffffc0000000, 80'h0000001ffffff8000000, 80'h000000ffc003ff000000, 80'h000003fc08703fc00000,
    80'h00000fe03cf807f00000, 80'h00003f003c1800fc0000, 80'h00007e000c18007f0000, 80'h0001f8000c38001f8000,
    80'h0003e0000c700007c000, 80'h0007c0000ce00003e000, 80'h000f00003ef80000f000, 80'h001e0000000000007800,
    80'h003c0000000000003c00, 80'h00780000000000001e00, 80'h00f00000000000000f00, 80'h01e00000000000000780,
    80'h01c000000000000003c0, 80'h03c000000000000003c0, 80'h078000000000000001e0, 80'h070000000000000000e0,
    80'h0f0000000000000000f0, 80'h0e000000000000000070, 80'h1e000000000000000038, 80'h1c00000000000000003c,
    80'h3800000000000000001c, 80'h3800000000000000001c, 80'h3800000000000000001e, 80'h7000000000000000000e,
    80'h7000000000000000000e, 80'h7000000000000000000e, 80'he0000000000000000007, 80'he0000000000000000007,
    80'he0000000000000000007, 80'he0000000000000000007, 80'hc0000000000000000003, 80'hc0000000000000000003,
    80'hc7000000000000000073, 80'hcf8000000000000000fb, 80'hcd80000000000000001b, 80'hcdc0000000000000003b,
    80'hcfc0000000000000007b, 80'hc780000000000000001b, 80'hc180000000000000009b, 80'hcf0000000000000000fb,
    80'hc0000000000000000003, 80'hc0000000000000000003, 80'he0000000000000000007, 80'he0000000000000000007,
    80'he0000000000000000007, 80'he0000000000000000007, 80'h7000000000000000000e, 80'h7000000000000000000e,
    80'h7000000000000000000e, 80'h3800000000000000001e, 80'h3800000000000000001c, 80'h3800000000000000001c,
    80'h1c00000000000000003c, 80'h1e000000000000000038, 80'h0e000000000000000070, 80'h0f0000000000000000f0,
    80'h070000000000000000e0, 80'h078000000000000001e0, 80'h03c000000000000001c0, 80'h03c000000000000003c0,
    80'h01e00000000000000780, 80'h00f00000000000000f00, 80'h00780000000000001e00, 80'h003c0000000000003c00,
    80'h001e0000000000007800, 80'h000f000000e00000f000, 80'h0007c00003e00001e000, 80'h0003e00003000007c000,
    80'h0001f80003e0001f8000, 80'h0000fc000370003f0000, 80'h00003f00037000fc0000, 80'h00000fe0036007f00000,
    80'h000003fc03e03fc00000, 80'h000001ffc003ff800000, 80'h0000003ffffffc000000, 80'h00000003ffffc0000000
};

wire [0:15] B_char [0:15] = '{
    16'h0000, 16'h0000, 16'h0000, 16'h3FF0, 16'h181C, 16'h180C, 16'h181C, 16'h1870,
    16'h1FB8, 16'h180C, 16'h180E, 16'h180E, 16'h180C, 16'hFFF0, 16'h0000, 16'h0000
};

wire [0:15] J_char [0:15] = '{
    16'h0000, 16'h0000, 16'h03FC, 16'h0060, 16'h0060, 16'h0060, 16'h0060, 16'h0060,
    16'h0060, 16'h0060, 16'h0060, 16'h0060, 16'h0060, 16'h70C0, 16'h1F00, 16'h0000
};

wire [0:15] S_char [0:15] = '{
    16'h0000, 16'h0000, 16'h0FF8, 16'h3008, 16'h2000, 16'h3000, 16'h1E00, 16'h01E0,
    16'h0018, 16'h000C, 16'h200C, 16'h3008, 16'h2FF0, 16'h0000, 16'h0000, 16'h0000
};

wire [0:15] N_char [0:15] = '{
    16'h0000, 16'h0000, 16'h780E, 16'h3C04, 16'h2E04, 16'h2704, 16'h2384, 16'h20C4,
    16'h2064, 16'h2034, 16'h201C, 16'h200C, 16'hF804, 16'h0000, 16'h0000, 16'h0000
};

wire [0:15] Y_char [0:15] = '{
    16'h0000, 16'h0000, 16'h381C, 16'h1808, 16'h0C10, 16'h0C20, 16'h0640, 16'h0340,
    16'h0180, 16'h0180, 16'h0180, 16'h0180, 16'h07E0, 16'h0000, 16'h0000, 16'h0000
};

wire [0:15] C_char [0:15] = '{
    16'h0000, 16'h0000, 16'h07FC, 16'h1804, 16'h3002, 16'h7000, 16'h6000, 16'h6000,
    16'h6000, 16'h7000, 16'h3002, 16'h180C, 16'h07F0, 16'h0000, 16'h0000, 16'h0000
};



    function automatic [15:0] get_minute_pixel;
        input [5:0] minute;
        input [15:0] x_pos;
        input [15:0] y_pos;
        begin
            case(minute)
                6'd0: get_minute_pixel = minute_000[y_pos][x_pos];
                6'd1: get_minute_pixel = minute_006[y_pos][x_pos];
                6'd2: get_minute_pixel = minute_012[y_pos][x_pos];
                6'd3: get_minute_pixel = minute_018[y_pos][x_pos];
                6'd4: get_minute_pixel = minute_024[y_pos][x_pos];
                6'd5: get_minute_pixel = minute_030[y_pos][x_pos];
                6'd6: get_minute_pixel = minute_036[y_pos][x_pos];
                6'd7: get_minute_pixel = minute_042[y_pos][x_pos];
                6'd8: get_minute_pixel = minute_048[y_pos][x_pos];
                6'd9: get_minute_pixel = minute_054[y_pos][x_pos];
                6'd10: get_minute_pixel = minute_060[y_pos][x_pos];
                6'd11: get_minute_pixel = minute_066[y_pos][x_pos];
                6'd12: get_minute_pixel = minute_072[y_pos][x_pos];
                6'd13: get_minute_pixel = minute_078[y_pos][x_pos];
                6'd14: get_minute_pixel = minute_084[y_pos][x_pos];
                6'd15: get_minute_pixel = minute_090[y_pos][x_pos];
                6'd16: get_minute_pixel = minute_096[y_pos][x_pos];
                6'd17: get_minute_pixel = minute_102[y_pos][x_pos];
                6'd18: get_minute_pixel = minute_108[y_pos][x_pos];
                6'd19: get_minute_pixel = minute_114[y_pos][x_pos];
                6'd20: get_minute_pixel = minute_120[y_pos][x_pos];
                6'd21: get_minute_pixel = minute_126[y_pos][x_pos];
                6'd22: get_minute_pixel = minute_132[y_pos][x_pos];
                6'd23: get_minute_pixel = minute_138[y_pos][x_pos];
                6'd24: get_minute_pixel = minute_144[y_pos][x_pos];
                6'd25: get_minute_pixel = minute_150[y_pos][x_pos];
                6'd26: get_minute_pixel = minute_156[y_pos][x_pos];
                6'd27: get_minute_pixel = minute_162[y_pos][x_pos];
                6'd28: get_minute_pixel = minute_168[y_pos][x_pos];
                6'd29: get_minute_pixel = minute_174[y_pos][x_pos];
                6'd30: get_minute_pixel = minute_180[y_pos][x_pos];
                6'd31: get_minute_pixel = minute_186[y_pos][x_pos];
                6'd32: get_minute_pixel = minute_192[y_pos][x_pos];
                6'd33: get_minute_pixel = minute_198[y_pos][x_pos];
                6'd34: get_minute_pixel = minute_204[y_pos][x_pos];
                6'd35: get_minute_pixel = minute_210[y_pos][x_pos];
                6'd36: get_minute_pixel = minute_216[y_pos][x_pos];
                6'd37: get_minute_pixel = minute_222[y_pos][x_pos];
                6'd38: get_minute_pixel = minute_228[y_pos][x_pos];
                6'd39: get_minute_pixel = minute_234[y_pos][x_pos];
                6'd40: get_minute_pixel = minute_240[y_pos][x_pos];
                6'd41: get_minute_pixel = minute_246[y_pos][x_pos];
                6'd42: get_minute_pixel = minute_252[y_pos][x_pos];
                6'd43: get_minute_pixel = minute_258[y_pos][x_pos];
                6'd44: get_minute_pixel = minute_264[y_pos][x_pos];
                6'd45: get_minute_pixel = minute_270[y_pos][x_pos];
                6'd46: get_minute_pixel = minute_276[y_pos][x_pos];
                6'd47: get_minute_pixel = minute_282[y_pos][x_pos];
                6'd48: get_minute_pixel = minute_288[y_pos][x_pos];
                6'd49: get_minute_pixel = minute_294[y_pos][x_pos];
                6'd50: get_minute_pixel = minute_300[y_pos][x_pos];
                6'd51: get_minute_pixel = minute_306[y_pos][x_pos];
                6'd52: get_minute_pixel = minute_312[y_pos][x_pos];
                6'd53: get_minute_pixel = minute_318[y_pos][x_pos];
                6'd54: get_minute_pixel = minute_324[y_pos][x_pos];
                6'd55: get_minute_pixel = minute_330[y_pos][x_pos];
                6'd56: get_minute_pixel = minute_336[y_pos][x_pos];
                6'd57: get_minute_pixel = minute_342[y_pos][x_pos];
                6'd58: get_minute_pixel = minute_348[y_pos][x_pos];
                6'd59: get_minute_pixel = minute_354[y_pos][x_pos];
                default: get_minute_pixel = 1'b0;
            endcase
        end
    endfunction

    function automatic [15:0] get_second_pixel;
        input [5:0] second;
        input [15:0] x_pos;
        input [15:0] y_pos;
        begin
            case(second)
                6'd0: get_second_pixel = second_000[y_pos][x_pos];
                6'd1: get_second_pixel = second_006[y_pos][x_pos];
                6'd2: get_second_pixel = second_012[y_pos][x_pos];
                6'd3: get_second_pixel = second_018[y_pos][x_pos];
                6'd4: get_second_pixel = second_024[y_pos][x_pos];
                6'd5: get_second_pixel = second_030[y_pos][x_pos];
                6'd6: get_second_pixel = second_036[y_pos][x_pos];
                6'd7: get_second_pixel = second_042[y_pos][x_pos];
                6'd8: get_second_pixel = second_048[y_pos][x_pos];
                6'd9: get_second_pixel = second_054[y_pos][x_pos];
                6'd10: get_second_pixel = second_060[y_pos][x_pos];
                6'd11: get_second_pixel = second_066[y_pos][x_pos];
                6'd12: get_second_pixel = second_072[y_pos][x_pos];
                6'd13: get_second_pixel = second_078[y_pos][x_pos];
                6'd14: get_second_pixel = second_084[y_pos][x_pos];
                6'd15: get_second_pixel = second_090[y_pos][x_pos];
                6'd16: get_second_pixel = second_096[y_pos][x_pos];
                6'd17: get_second_pixel = second_102[y_pos][x_pos];
                6'd18: get_second_pixel = second_108[y_pos][x_pos];
                6'd19: get_second_pixel = second_114[y_pos][x_pos];
                6'd20: get_second_pixel = second_120[y_pos][x_pos];
                6'd21: get_second_pixel = second_126[y_pos][x_pos];
                6'd22: get_second_pixel = second_132[y_pos][x_pos];
                6'd23: get_second_pixel = second_138[y_pos][x_pos];
                6'd24: get_second_pixel = second_144[y_pos][x_pos];
                6'd25: get_second_pixel = second_150[y_pos][x_pos];
                6'd26: get_second_pixel = second_156[y_pos][x_pos];
                6'd27: get_second_pixel = second_162[y_pos][x_pos];
                6'd28: get_second_pixel = second_168[y_pos][x_pos];
                6'd29: get_second_pixel = second_174[y_pos][x_pos];
                6'd30: get_second_pixel = second_180[y_pos][x_pos];
                6'd31: get_second_pixel = second_186[y_pos][x_pos];
                6'd32: get_second_pixel = second_192[y_pos][x_pos];
                6'd33: get_second_pixel = second_198[y_pos][x_pos];
                6'd34: get_second_pixel = second_204[y_pos][x_pos];
                6'd35: get_second_pixel = second_210[y_pos][x_pos];
                6'd36: get_second_pixel = second_216[y_pos][x_pos];
                6'd37: get_second_pixel = second_222[y_pos][x_pos];
                6'd38: get_second_pixel = second_228[y_pos][x_pos];
                6'd39: get_second_pixel = second_234[y_pos][x_pos];
                6'd40: get_second_pixel = second_240[y_pos][x_pos];
                6'd41: get_second_pixel = second_246[y_pos][x_pos];
                6'd42: get_second_pixel = second_252[y_pos][x_pos];
                6'd43: get_second_pixel = second_258[y_pos][x_pos];
                6'd44: get_second_pixel = second_264[y_pos][x_pos];
                6'd45: get_second_pixel = second_270[y_pos][x_pos];
                6'd46: get_second_pixel = second_276[y_pos][x_pos];
                6'd47: get_second_pixel = second_282[y_pos][x_pos];
                6'd48: get_second_pixel = second_288[y_pos][x_pos];
                6'd49: get_second_pixel = second_294[y_pos][x_pos];
                6'd50: get_second_pixel = second_300[y_pos][x_pos];
                6'd51: get_second_pixel = second_306[y_pos][x_pos];
                6'd52: get_second_pixel = second_312[y_pos][x_pos];
                6'd53: get_second_pixel = second_318[y_pos][x_pos];
                6'd54: get_second_pixel = second_324[y_pos][x_pos];
                6'd55: get_second_pixel = second_330[y_pos][x_pos];
                6'd56: get_second_pixel = second_336[y_pos][x_pos];
                6'd57: get_second_pixel = second_342[y_pos][x_pos];
                6'd58: get_second_pixel = second_348[y_pos][x_pos];
                6'd59: get_second_pixel = second_354[y_pos][x_pos];
                default: get_second_pixel = 1'b0;
            endcase
        end
    endfunction

    function automatic [15:0] get_hour_pixel;
        input [5:0] hour;
        input [15:0] x_pos;
        input [15:0] y_pos;
        begin
            case(hour)
                6'd0: get_hour_pixel = hour_000[y_pos][x_pos];
                6'd1: get_hour_pixel = hour_030[y_pos][x_pos];
                6'd2: get_hour_pixel = hour_060[y_pos][x_pos];
                6'd3: get_hour_pixel = hour_090[y_pos][x_pos];
                6'd4: get_hour_pixel = hour_120[y_pos][x_pos];
                6'd5: get_hour_pixel = hour_150[y_pos][x_pos];
                6'd6: get_hour_pixel = hour_180[y_pos][x_pos];
                6'd7: get_hour_pixel = hour_210[y_pos][x_pos];
                6'd8: get_hour_pixel = hour_240[y_pos][x_pos];
                6'd9: get_hour_pixel = hour_270[y_pos][x_pos];
                6'd10: get_hour_pixel = hour_300[y_pos][x_pos];
                6'd11: get_hour_pixel = hour_330[y_pos][x_pos];
      
                default: get_hour_pixel = 1'b0;
            endcase
        end
    endfunction

always @(posedge PixelClk or negedge nRST) begin
    if(!nRST) begin
        LCD_R <= 5'b11111;
        LCD_G <= 6'b111111;
        LCD_B <= 5'b11111;
    end
    else begin




        if(PixelCount >= 600 && PixelCount < 680 && LineCount >= 180 && LineCount < 260) begin
            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 600;
            y_pos = LineCount - 180;
            
           // 默认背景色
            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;
            
            if(clock[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end

          // 时针
            if(get_hour_pixel(hour_decimal%12, x_pos, y_pos)) begin
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b11111;
            end


            // 分针
            if(get_minute_pixel(minute_decimal, x_pos, y_pos)) begin
                LCD_R <= 5'b00000;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b00000;
            end
            
            // 再检查秒针，这样秒针会覆盖分针
            if(get_second_pixel(second_decimal, x_pos, y_pos)) begin 
                LCD_R <= 5'b11111;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
        end


        else if(PixelCount >= 780 && PixelCount < 860 && LineCount >= 180 && LineCount < 260) begin 
            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 780;
            y_pos = LineCount - 180;
            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;


            if(clock[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end

            if(get_hour_pixel((hour_decimal-12)%12, x_pos, y_pos)) begin
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b11111;
            end

            if(get_minute_pixel((minute_decimal)%60, x_pos, y_pos)) begin
                LCD_R <= 5'b00000;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b00000;
            end

            if(get_second_pixel((second_decimal)%60, x_pos, y_pos)) begin 
                LCD_R <= 5'b11111;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
        
        end

        else if(PixelCount >= 610 && PixelCount < 626 && LineCount >= 270 && LineCount < 286) begin

            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 610;
            y_pos = LineCount - 270;

            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;

            if(B_char[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end
        end

        else if(PixelCount >= 630 && PixelCount < 646 && LineCount >= 270 && LineCount < 286) begin

            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 630;
            y_pos = LineCount - 270;

            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;

            if(J_char[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end
        end

        else if(PixelCount >= 650 && PixelCount < 666 && LineCount >= 270 && LineCount < 286) begin

            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 650;
            y_pos = LineCount - 270;

            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;

            if(S_char[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end
        end
            

        else if(PixelCount >= 790 && PixelCount < 806 && LineCount >= 270 && LineCount < 286) begin

            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 790;
            y_pos = LineCount - 270;

            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;

            if(N_char[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end
        end

        else if(PixelCount >= 810 && PixelCount < 826 && LineCount >= 270 && LineCount < 286) begin

            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 810;
            y_pos = LineCount - 270;

            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;

            if(Y_char[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end
        end

        else if(PixelCount >= 830 && PixelCount < 846 && LineCount >= 270 && LineCount < 286) begin

            integer x_pos;
            integer y_pos;
            x_pos = PixelCount - 830;
            y_pos = LineCount - 270;

            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;

            if(C_char[y_pos][x_pos] == 1'b1) begin 
                LCD_R <= 5'b00000;
                LCD_G <= 6'b000000;
                LCD_B <= 5'b00000;
            end
            else begin
                LCD_R <= 5'b11111;
                LCD_G <= 6'b111111;
                LCD_B <= 5'b11111;
            end
        end


        else begin
            LCD_R <= 5'b11111;
            LCD_G <= 6'b111111;
            LCD_B <= 5'b11111;
        end
    end

end
endmodule